../../idram_xilinx.vhd