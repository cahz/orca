../../../rtl/components.vhd