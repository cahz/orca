../../bram_xilinx.vhd