../../../rtl/iram_microsemi.vhd