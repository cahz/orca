../../rtl/decode.vhd