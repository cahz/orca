../../rtl/orca_core.vhd