../../../rtl/cache_mux.vhd