../../../rtl/bram_xilinx.vhd