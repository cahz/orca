../../rtl/execute.vhd