../../../rtl/icache.vhd