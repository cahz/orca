../../../rtl/axi_instruction_master.vhd