../../rtl/alu.vhd