-- Version: 
-- VHDL Black Box file 
-- 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity MSS_120 is
	generic (
		INIT:std_logic_vector := x"0";
		ACT_UBITS:std_logic_vector := x"0";
		MEMORYFILE:string := "";
		RTC_MAIN_XTL_FREQ:real := 0.0;
		RTC_MAIN_XTL_MODE:string := "";
		DDR_CLK_FREQ:real := 0.0	);
   port( 
       CAN_RXBUS_MGPIO3A_H2F_A : out std_logic;
       CAN_RXBUS_MGPIO3A_H2F_B : out std_logic;
       CAN_TX_EBL_MGPIO4A_H2F_A : out std_logic;
       CAN_TX_EBL_MGPIO4A_H2F_B : out std_logic;
       CAN_TXBUS_MGPIO2A_H2F_A : out std_logic;
       CAN_TXBUS_MGPIO2A_H2F_B : out std_logic;
       CLK_CONFIG_APB : out std_logic;
       COMMS_INT : out std_logic;
       CONFIG_PRESET_N : out std_logic;
       EDAC_ERROR : out std_logic_vector(7 downto 0);
       F_FM0_RDATA : out std_logic_vector(31 downto 0);
       F_FM0_READYOUT : out std_logic;
       F_FM0_RESP : out std_logic;
       F_FM1_RDATA : out std_logic_vector(31 downto 0);
       F_FM1_READYOUT : out std_logic;
       F_FM1_RESP : out std_logic;
       F_HM0_ADDR : out std_logic_vector(31 downto 0);
       F_HM0_ENABLE : out std_logic;
       F_HM0_SEL : out std_logic;
       F_HM0_SIZE : out std_logic_vector(1 downto 0);
       F_HM0_TRANS1 : out std_logic;
       F_HM0_WDATA : out std_logic_vector(31 downto 0);
       F_HM0_WRITE : out std_logic;
       F_HM1_ADDR : out std_logic_vector(31 downto 0);
       F_HM1_ENABLE : out std_logic;
       F_HM1_SEL : out std_logic;
       F_HM1_SIZE : out std_logic_vector(1 downto 0);
       F_HM1_TRANS1 : out std_logic;
       F_HM1_WDATA : out std_logic_vector(31 downto 0);
       F_HM1_WRITE : out std_logic;
       FAB_CHRGVBUS : out std_logic;
       FAB_DISCHRGVBUS : out std_logic;
       FAB_DMPULLDOWN : out std_logic;
       FAB_DPPULLDOWN : out std_logic;
       FAB_DRVVBUS : out std_logic;
       FAB_IDPULLUP : out std_logic;
       FAB_OPMODE : out std_logic_vector(1 downto 0);
       FAB_SUSPENDM : out std_logic;
       FAB_TERMSEL : out std_logic;
       FAB_TXVALID : out std_logic;
       FAB_VCONTROL : out std_logic_vector(3 downto 0);
       FAB_VCONTROLLOADM : out std_logic;
       FAB_XCVRSEL : out std_logic_vector(1 downto 0);
       FAB_XDATAOUT : out std_logic_vector(7 downto 0);
       FACC_GLMUX_SEL : out std_logic;
       FIC32_0_MASTER : out std_logic_vector(1 downto 0);
       FIC32_1_MASTER : out std_logic_vector(1 downto 0);
       FPGA_RESET_N : out std_logic;
       GTX_CLK : out std_logic;
       H2F_INTERRUPT : out std_logic_vector(15 downto 0);
       H2F_NMI : out std_logic;
       H2FCALIB : out std_logic;
       I2C0_SCL_MGPIO31B_H2F_A : out std_logic;
       I2C0_SCL_MGPIO31B_H2F_B : out std_logic;
       I2C0_SDA_MGPIO30B_H2F_A : out std_logic;
       I2C0_SDA_MGPIO30B_H2F_B : out std_logic;
       I2C1_SCL_MGPIO1A_H2F_A : out std_logic;
       I2C1_SCL_MGPIO1A_H2F_B : out std_logic;
       I2C1_SDA_MGPIO0A_H2F_A : out std_logic;
       I2C1_SDA_MGPIO0A_H2F_B : out std_logic;
       MDCF : out std_logic;
       MDOENF : out std_logic;
       MDOF : out std_logic;
       MMUART0_CTS_MGPIO19B_H2F_A : out std_logic;
       MMUART0_CTS_MGPIO19B_H2F_B : out std_logic;
       MMUART0_DCD_MGPIO22B_H2F_A : out std_logic;
       MMUART0_DCD_MGPIO22B_H2F_B : out std_logic;
       MMUART0_DSR_MGPIO20B_H2F_A : out std_logic;
       MMUART0_DSR_MGPIO20B_H2F_B : out std_logic;
       MMUART0_DTR_MGPIO18B_H2F_A : out std_logic;
       MMUART0_DTR_MGPIO18B_H2F_B : out std_logic;
       MMUART0_RI_MGPIO21B_H2F_A : out std_logic;
       MMUART0_RI_MGPIO21B_H2F_B : out std_logic;
       MMUART0_RTS_MGPIO17B_H2F_A : out std_logic;
       MMUART0_RTS_MGPIO17B_H2F_B : out std_logic;
       MMUART0_RXD_MGPIO28B_H2F_A : out std_logic;
       MMUART0_RXD_MGPIO28B_H2F_B : out std_logic;
       MMUART0_SCK_MGPIO29B_H2F_A : out std_logic;
       MMUART0_SCK_MGPIO29B_H2F_B : out std_logic;
       MMUART0_TXD_MGPIO27B_H2F_A : out std_logic;
       MMUART0_TXD_MGPIO27B_H2F_B : out std_logic;
       MMUART1_DTR_MGPIO12B_H2F_A : out std_logic;
       MMUART1_RTS_MGPIO11B_H2F_A : out std_logic;
       MMUART1_RTS_MGPIO11B_H2F_B : out std_logic;
       MMUART1_RXD_MGPIO26B_H2F_A : out std_logic;
       MMUART1_RXD_MGPIO26B_H2F_B : out std_logic;
       MMUART1_SCK_MGPIO25B_H2F_A : out std_logic;
       MMUART1_SCK_MGPIO25B_H2F_B : out std_logic;
       MMUART1_TXD_MGPIO24B_H2F_A : out std_logic;
       MMUART1_TXD_MGPIO24B_H2F_B : out std_logic;
       MPLL_LOCK : out std_logic;
       PER2_FABRIC_PADDR : out std_logic_vector(16 downto 2);
       PER2_FABRIC_PENABLE : out std_logic;
       PER2_FABRIC_PSEL : out std_logic;
       PER2_FABRIC_PWDATA : out std_logic_vector(31 downto 0);
       PER2_FABRIC_PWRITE : out std_logic;
       RTC_MATCH : out std_logic;
       SLEEPDEEP : out std_logic;
       SLEEPHOLDACK : out std_logic;
       SLEEPING : out std_logic;
       SMBALERT_NO0 : out std_logic;
       SMBALERT_NO1 : out std_logic;
       SMBSUS_NO0 : out std_logic;
       SMBSUS_NO1 : out std_logic;
       SPI0_CLK_OUT : out std_logic;
       SPI0_SDI_MGPIO5A_H2F_A : out std_logic;
       SPI0_SDI_MGPIO5A_H2F_B : out std_logic;
       SPI0_SDO_MGPIO6A_H2F_A : out std_logic;
       SPI0_SDO_MGPIO6A_H2F_B : out std_logic;
       SPI0_SS0_MGPIO7A_H2F_A : out std_logic;
       SPI0_SS0_MGPIO7A_H2F_B : out std_logic;
       SPI0_SS1_MGPIO8A_H2F_A : out std_logic;
       SPI0_SS1_MGPIO8A_H2F_B : out std_logic;
       SPI0_SS2_MGPIO9A_H2F_A : out std_logic;
       SPI0_SS2_MGPIO9A_H2F_B : out std_logic;
       SPI0_SS3_MGPIO10A_H2F_A : out std_logic;
       SPI0_SS3_MGPIO10A_H2F_B : out std_logic;
       SPI0_SS4_MGPIO19A_H2F_A : out std_logic;
       SPI0_SS5_MGPIO20A_H2F_A : out std_logic;
       SPI0_SS6_MGPIO21A_H2F_A : out std_logic;
       SPI0_SS7_MGPIO22A_H2F_A : out std_logic;
       SPI1_CLK_OUT : out std_logic;
       SPI1_SDI_MGPIO11A_H2F_A : out std_logic;
       SPI1_SDI_MGPIO11A_H2F_B : out std_logic;
       SPI1_SDO_MGPIO12A_H2F_A : out std_logic;
       SPI1_SDO_MGPIO12A_H2F_B : out std_logic;
       SPI1_SS0_MGPIO13A_H2F_A : out std_logic;
       SPI1_SS0_MGPIO13A_H2F_B : out std_logic;
       SPI1_SS1_MGPIO14A_H2F_A : out std_logic;
       SPI1_SS1_MGPIO14A_H2F_B : out std_logic;
       SPI1_SS2_MGPIO15A_H2F_A : out std_logic;
       SPI1_SS2_MGPIO15A_H2F_B : out std_logic;
       SPI1_SS3_MGPIO16A_H2F_A : out std_logic;
       SPI1_SS3_MGPIO16A_H2F_B : out std_logic;
       SPI1_SS4_MGPIO17A_H2F_A : out std_logic;
       SPI1_SS5_MGPIO18A_H2F_A : out std_logic;
       SPI1_SS6_MGPIO23A_H2F_A : out std_logic;
       SPI1_SS7_MGPIO24A_H2F_A : out std_logic;
       TCGF : out std_logic_vector(9 downto 0);
       TRACECLK : out std_logic;
       TRACEDATA : out std_logic_vector(3 downto 0);
       TX_CLK : out std_logic;
       TX_ENF : out std_logic;
       TX_ERRF : out std_logic;
       TXCTL_EN_RIF : out std_logic;
       TXD_RIF : out std_logic_vector(3 downto 0);
       TXDF : out std_logic_vector(7 downto 0);
       TXEV : out std_logic;
       WDOGTIMEOUT : out std_logic;
       F_ARREADY_HREADYOUT1 : out std_logic;
       F_AWREADY_HREADYOUT0 : out std_logic;
       F_BID : out std_logic_vector(3 downto 0);
       F_BRESP_HRESP0 : out std_logic_vector(1 downto 0);
       F_BVALID : out std_logic;
       F_RDATA_HRDATA01 : out std_logic_vector(63 downto 0);
       F_RID : out std_logic_vector(3 downto 0);
       F_RLAST : out std_logic;
       F_RRESP_HRESP1 : out std_logic_vector(1 downto 0);
       F_RVALID : out std_logic;
       F_WREADY : out std_logic;
       MDDR_FABRIC_PRDATA : out std_logic_vector(15 downto 0);
       MDDR_FABRIC_PREADY : out std_logic;
       MDDR_FABRIC_PSLVERR : out std_logic;
       REV_ARADDR : out std_logic_vector(31 downto 0);
       REV_ARBURST : out std_logic_vector(1 downto 0);
       REV_ARID : out std_logic_vector(3 downto 0);
       REV_ARLEN : out std_logic_vector(3 downto 0);
       REV_ARLOCK : out std_logic_vector(1 downto 0);
       REV_ARSIZE : out std_logic_vector(1 downto 0);
       REV_AWADDR : out std_logic_vector(31 downto 0);
       REV_AWLOCK : out std_logic_vector(1 downto 0);
       REV_AWSIZE : out std_logic_vector(1 downto 0);
       REV_RREADY : out std_logic;
       REV_WID : out std_logic_vector(3 downto 0);
       REV_WSTRB : out std_logic_vector(7 downto 0);
       CAN_RXBUS_F2H_SCP : in std_logic;
       CAN_TX_EBL_F2H_SCP : in std_logic;
       CAN_TXBUS_F2H_SCP : in std_logic;
       CLK_BASE : in std_logic;
       COLF : in std_logic;
       CRSF : in std_logic;
       F2_DMAREADY : in std_logic_vector(1 downto 0);
       F2H_INTERRUPT : in std_logic_vector(15 downto 0);
       F2HCALIB : in std_logic;
       F_DMAREADY : in std_logic_vector(1 downto 0);
       F_FM0_ADDR : in std_logic_vector(31 downto 0);
       F_FM0_ENABLE : in std_logic;
       F_FM0_MASTLOCK : in std_logic;
       F_FM0_READY : in std_logic;
       F_FM0_SEL : in std_logic;
       F_FM0_SIZE : in std_logic_vector(1 downto 0);
       F_FM0_TRANS1 : in std_logic;
       F_FM0_WDATA : in std_logic_vector(31 downto 0);
       F_FM0_WRITE : in std_logic;
       F_FM1_ADDR : in std_logic_vector(31 downto 0);
       F_FM1_ENABLE : in std_logic;
       F_FM1_MASTLOCK : in std_logic;
       F_FM1_READY : in std_logic;
       F_FM1_SEL : in std_logic;
       F_FM1_SIZE : in std_logic_vector(1 downto 0);
       F_FM1_TRANS1 : in std_logic;
       F_FM1_WDATA : in std_logic_vector(31 downto 0);
       F_FM1_WRITE : in std_logic;
       F_HM0_RDATA : in std_logic_vector(31 downto 0);
       F_HM0_READY : in std_logic;
       F_HM0_RESP : in std_logic;
       F_HM1_RDATA : in std_logic_vector(31 downto 0);
       F_HM1_READY : in std_logic;
       F_HM1_RESP : in std_logic;
       FAB_AVALID : in std_logic;
       FAB_HOSTDISCON : in std_logic;
       FAB_IDDIG : in std_logic;
       FAB_LINESTATE : in std_logic_vector(1 downto 0);
       FAB_M3_RESET_N : in std_logic;
       FAB_PLL_LOCK : in std_logic;
       FAB_RXACTIVE : in std_logic;
       FAB_RXERROR : in std_logic;
       FAB_RXVALID : in std_logic;
       FAB_RXVALIDH : in std_logic;
       FAB_SESSEND : in std_logic;
       FAB_TXREADY : in std_logic;
       FAB_VBUSVALID : in std_logic;
       FAB_VSTATUS : in std_logic_vector(7 downto 0);
       FAB_XDATAIN : in std_logic_vector(7 downto 0);
       GTX_CLKPF : in std_logic;
       I2C0_BCLK : in std_logic;
       I2C0_SCL_F2H_SCP : in std_logic;
       I2C0_SDA_F2H_SCP : in std_logic;
       I2C1_BCLK : in std_logic;
       I2C1_SCL_F2H_SCP : in std_logic;
       I2C1_SDA_F2H_SCP : in std_logic;
       MDIF : in std_logic;
       MGPIO0A_F2H_GPIN : in std_logic;
       MGPIO10A_F2H_GPIN : in std_logic;
       MGPIO11A_F2H_GPIN : in std_logic;
       MGPIO11B_F2H_GPIN : in std_logic;
       MGPIO12A_F2H_GPIN : in std_logic;
       MGPIO13A_F2H_GPIN : in std_logic;
       MGPIO14A_F2H_GPIN : in std_logic;
       MGPIO15A_F2H_GPIN : in std_logic;
       MGPIO16A_F2H_GPIN : in std_logic;
       MGPIO17B_F2H_GPIN : in std_logic;
       MGPIO18B_F2H_GPIN : in std_logic;
       MGPIO19B_F2H_GPIN : in std_logic;
       MGPIO1A_F2H_GPIN : in std_logic;
       MGPIO20B_F2H_GPIN : in std_logic;
       MGPIO21B_F2H_GPIN : in std_logic;
       MGPIO22B_F2H_GPIN : in std_logic;
       MGPIO24B_F2H_GPIN : in std_logic;
       MGPIO25B_F2H_GPIN : in std_logic;
       MGPIO26B_F2H_GPIN : in std_logic;
       MGPIO27B_F2H_GPIN : in std_logic;
       MGPIO28B_F2H_GPIN : in std_logic;
       MGPIO29B_F2H_GPIN : in std_logic;
       MGPIO2A_F2H_GPIN : in std_logic;
       MGPIO30B_F2H_GPIN : in std_logic;
       MGPIO31B_F2H_GPIN : in std_logic;
       MGPIO3A_F2H_GPIN : in std_logic;
       MGPIO4A_F2H_GPIN : in std_logic;
       MGPIO5A_F2H_GPIN : in std_logic;
       MGPIO6A_F2H_GPIN : in std_logic;
       MGPIO7A_F2H_GPIN : in std_logic;
       MGPIO8A_F2H_GPIN : in std_logic;
       MGPIO9A_F2H_GPIN : in std_logic;
       MMUART0_CTS_F2H_SCP : in std_logic;
       MMUART0_DCD_F2H_SCP : in std_logic;
       MMUART0_DSR_F2H_SCP : in std_logic;
       MMUART0_DTR_F2H_SCP : in std_logic;
       MMUART0_RI_F2H_SCP : in std_logic;
       MMUART0_RTS_F2H_SCP : in std_logic;
       MMUART0_RXD_F2H_SCP : in std_logic;
       MMUART0_SCK_F2H_SCP : in std_logic;
       MMUART0_TXD_F2H_SCP : in std_logic;
       MMUART1_CTS_F2H_SCP : in std_logic;
       MMUART1_DCD_F2H_SCP : in std_logic;
       MMUART1_DSR_F2H_SCP : in std_logic;
       MMUART1_RI_F2H_SCP : in std_logic;
       MMUART1_RTS_F2H_SCP : in std_logic;
       MMUART1_RXD_F2H_SCP : in std_logic;
       MMUART1_SCK_F2H_SCP : in std_logic;
       MMUART1_TXD_F2H_SCP : in std_logic;
       PER2_FABRIC_PRDATA : in std_logic_vector(31 downto 0);
       PER2_FABRIC_PREADY : in std_logic;
       PER2_FABRIC_PSLVERR : in std_logic;
       RCGF : in std_logic_vector(9 downto 0);
       RX_CLKPF : in std_logic;
       RX_DVF : in std_logic;
       RX_ERRF : in std_logic;
       RX_EV : in std_logic;
       RXDF : in std_logic_vector(7 downto 0);
       SLEEPHOLDREQ : in std_logic;
       SMBALERT_NI0 : in std_logic;
       SMBALERT_NI1 : in std_logic;
       SMBSUS_NI0 : in std_logic;
       SMBSUS_NI1 : in std_logic;
       SPI0_CLK_IN : in std_logic;
       SPI0_SDI_F2H_SCP : in std_logic;
       SPI0_SDO_F2H_SCP : in std_logic;
       SPI0_SS0_F2H_SCP : in std_logic;
       SPI0_SS1_F2H_SCP : in std_logic;
       SPI0_SS2_F2H_SCP : in std_logic;
       SPI0_SS3_F2H_SCP : in std_logic;
       SPI1_CLK_IN : in std_logic;
       SPI1_SDI_F2H_SCP : in std_logic;
       SPI1_SDO_F2H_SCP : in std_logic;
       SPI1_SS0_F2H_SCP : in std_logic;
       SPI1_SS1_F2H_SCP : in std_logic;
       SPI1_SS2_F2H_SCP : in std_logic;
       SPI1_SS3_F2H_SCP : in std_logic;
       TX_CLKPF : in std_logic;
       USER_MSS_GPIO_RESET_N : in std_logic;
       USER_MSS_RESET_N : in std_logic;
       XCLK_FAB : in std_logic;
       CLK_MDDR_APB : in std_logic;
       F_ARADDR_HADDR1 : in std_logic_vector(31 downto 0);
       F_ARBURST_HTRANS1 : in std_logic_vector(1 downto 0);
       F_ARID_HSEL1 : in std_logic_vector(3 downto 0);
       F_ARLEN_HBURST1 : in std_logic_vector(3 downto 0);
       F_ARLOCK_HMASTLOCK1 : in std_logic_vector(1 downto 0);
       F_ARSIZE_HSIZE1 : in std_logic_vector(1 downto 0);
       F_ARVALID_HWRITE1 : in std_logic;
       F_AWADDR_HADDR0 : in std_logic_vector(31 downto 0);
       F_AWBURST_HTRANS0 : in std_logic_vector(1 downto 0);
       F_AWID_HSEL0 : in std_logic_vector(3 downto 0);
       F_AWLEN_HBURST0 : in std_logic_vector(3 downto 0);
       F_AWLOCK_HMASTLOCK0 : in std_logic_vector(1 downto 0);
       F_AWSIZE_HSIZE0 : in std_logic_vector(1 downto 0);
       F_AWVALID_HWRITE0 : in std_logic;
       F_BREADY : in std_logic;
       F_RMW_AXI : in std_logic;
       F_RREADY : in std_logic;
       F_WDATA_HWDATA01 : in std_logic_vector(63 downto 0);
       F_WID_HREADY01 : in std_logic_vector(3 downto 0);
       F_WLAST : in std_logic;
       F_WSTRB : in std_logic_vector(7 downto 0);
       F_WVALID : in std_logic;
       FPGA_MDDR_ARESET_N : in std_logic;
       MDDR_FABRIC_PADDR : in std_logic_vector(10 downto 2);
       MDDR_FABRIC_PENABLE : in std_logic;
       MDDR_FABRIC_PSEL : in std_logic;
       MDDR_FABRIC_PWDATA : in std_logic_vector(15 downto 0);
       MDDR_FABRIC_PWRITE : in std_logic;
       PRESET_N : in std_logic;
       CAN_RXBUS_USBA_DATA1_MGPIO3A_IN : in std_logic;
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN : in std_logic;
       CAN_TXBUS_USBA_DATA0_MGPIO2A_IN : in std_logic;
       DM_IN : in std_logic_vector(4 downto 0);
       DRAM_DQ_IN : in std_logic_vector(35 downto 0);
       DRAM_DQS_IN : in std_logic_vector(4 downto 0);
       DRAM_FIFO_WE_IN : in std_logic_vector(2 downto 0);
       I2C0_SCL_USBC_DATA1_MGPIO31B_IN : in std_logic;
       I2C0_SDA_USBC_DATA0_MGPIO30B_IN : in std_logic;
       I2C1_SCL_USBA_DATA4_MGPIO1A_IN : in std_logic;
       I2C1_SDA_USBA_DATA3_MGPIO0A_IN : in std_logic;
       MGPIO0B_IN : in std_logic;
       MGPIO10B_IN : in std_logic;
       MGPIO1B_IN : in std_logic;
       MGPIO25A_IN : in std_logic;
       MGPIO26A_IN : in std_logic;
       MGPIO27A_IN : in std_logic;
       MGPIO28A_IN : in std_logic;
       MGPIO29A_IN : in std_logic;
       MGPIO2B_IN : in std_logic;
       MGPIO30A_IN : in std_logic;
       MGPIO31A_IN : in std_logic;
       MGPIO3B_IN : in std_logic;
       MGPIO4B_IN : in std_logic;
       MGPIO5B_IN : in std_logic;
       MGPIO6B_IN : in std_logic;
       MGPIO7B_IN : in std_logic;
       MGPIO8B_IN : in std_logic;
       MGPIO9B_IN : in std_logic;
       MMUART0_CTS_USBC_DATA7_MGPIO19B_IN : in std_logic;
       MMUART0_DCD_MGPIO22B_IN : in std_logic;
       MMUART0_DSR_MGPIO20B_IN : in std_logic;
       MMUART0_DTR_USBC_DATA6_MGPIO18B_IN : in std_logic;
       MMUART0_RI_MGPIO21B_IN : in std_logic;
       MMUART0_RTS_USBC_DATA5_MGPIO17B_IN : in std_logic;
       MMUART0_RXD_USBC_STP_MGPIO28B_IN : in std_logic;
       MMUART0_SCK_USBC_NXT_MGPIO29B_IN : in std_logic;
       MMUART0_TXD_USBC_DIR_MGPIO27B_IN : in std_logic;
       MMUART1_CTS_MGPIO13B_IN : in std_logic;
       MMUART1_DCD_MGPIO16B_IN : in std_logic;
       MMUART1_DSR_MGPIO14B_IN : in std_logic;
       MMUART1_DTR_MGPIO12B_IN : in std_logic;
       MMUART1_RI_MGPIO15B_IN : in std_logic;
       MMUART1_RTS_MGPIO11B_IN : in std_logic;
       MMUART1_RXD_USBC_DATA3_MGPIO26B_IN : in std_logic;
       MMUART1_SCK_USBC_DATA4_MGPIO25B_IN : in std_logic;
       MMUART1_TXD_USBC_DATA2_MGPIO24B_IN : in std_logic;
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN : in std_logic;
       RGMII_MDC_RMII_MDC_IN : in std_logic;
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN : in std_logic;
       RGMII_RX_CLK_IN : in std_logic;
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN : in std_logic;
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN : in std_logic;
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN : in std_logic;
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN : in std_logic;
       RGMII_RXD3_USBB_DATA4_IN : in std_logic;
       RGMII_TX_CLK_IN : in std_logic;
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN : in std_logic;
       RGMII_TXD0_RMII_TXD0_USBB_DIR_IN : in std_logic;
       RGMII_TXD1_RMII_TXD1_USBB_STP_IN : in std_logic;
       RGMII_TXD2_USBB_DATA5_IN : in std_logic;
       RGMII_TXD3_USBB_DATA6_IN : in std_logic;
       SPI0_SCK_USBA_XCLK_IN : in std_logic;
       SPI0_SDI_USBA_DIR_MGPIO5A_IN : in std_logic;
       SPI0_SDO_USBA_STP_MGPIO6A_IN : in std_logic;
       SPI0_SS0_USBA_NXT_MGPIO7A_IN : in std_logic;
       SPI0_SS1_USBA_DATA5_MGPIO8A_IN : in std_logic;
       SPI0_SS2_USBA_DATA6_MGPIO9A_IN : in std_logic;
       SPI0_SS3_USBA_DATA7_MGPIO10A_IN : in std_logic;
       SPI0_SS4_MGPIO19A_IN : in std_logic;
       SPI0_SS5_MGPIO20A_IN : in std_logic;
       SPI0_SS6_MGPIO21A_IN : in std_logic;
       SPI0_SS7_MGPIO22A_IN : in std_logic;
       SPI1_SCK_IN : in std_logic;
       SPI1_SDI_MGPIO11A_IN : in std_logic;
       SPI1_SDO_MGPIO12A_IN : in std_logic;
       SPI1_SS0_MGPIO13A_IN : in std_logic;
       SPI1_SS1_MGPIO14A_IN : in std_logic;
       SPI1_SS2_MGPIO15A_IN : in std_logic;
       SPI1_SS3_MGPIO16A_IN : in std_logic;
       SPI1_SS4_MGPIO17A_IN : in std_logic;
       SPI1_SS5_MGPIO18A_IN : in std_logic;
       SPI1_SS6_MGPIO23A_IN : in std_logic;
       SPI1_SS7_MGPIO24A_IN : in std_logic;
       USBC_XCLK_IN : in std_logic;
       USBD_DATA0_IN : in std_logic;
       USBD_DATA1_IN : in std_logic;
       USBD_DATA2_IN : in std_logic;
       USBD_DATA3_IN : in std_logic;
       USBD_DATA4_IN : in std_logic;
       USBD_DATA5_IN : in std_logic;
       USBD_DATA6_IN : in std_logic;
       USBD_DATA7_MGPIO23B_IN : in std_logic;
       USBD_DIR_IN : in std_logic;
       USBD_NXT_IN : in std_logic;
       USBD_STP_IN : in std_logic;
       USBD_XCLK_IN : in std_logic;
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT : out std_logic;
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT : out std_logic;
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT : out std_logic;
       DRAM_ADDR : out std_logic_vector(15 downto 0);
       DRAM_BA : out std_logic_vector(2 downto 0);
       DRAM_CASN : out std_logic;
       DRAM_CKE : out std_logic;
       DRAM_CLK : out std_logic;
       DRAM_CSN : out std_logic;
       DRAM_DM_RDQS_OUT : out std_logic_vector(4 downto 0);
       DRAM_DQ_OUT : out std_logic_vector(35 downto 0);
       DRAM_DQS_OUT : out std_logic_vector(4 downto 0);
       DRAM_FIFO_WE_OUT : out std_logic_vector(2 downto 0);
       DRAM_ODT : out std_logic;
       DRAM_RASN : out std_logic;
       DRAM_RSTN : out std_logic;
       DRAM_WEN : out std_logic;
       I2C0_SCL_USBC_DATA1_MGPIO31B_OUT : out std_logic;
       I2C0_SDA_USBC_DATA0_MGPIO30B_OUT : out std_logic;
       I2C1_SCL_USBA_DATA4_MGPIO1A_OUT : out std_logic;
       I2C1_SDA_USBA_DATA3_MGPIO0A_OUT : out std_logic;
       MGPIO0B_OUT : out std_logic;
       MGPIO10B_OUT : out std_logic;
       MGPIO1B_OUT : out std_logic;
       MGPIO25A_OUT : out std_logic;
       MGPIO26A_OUT : out std_logic;
       MGPIO27A_OUT : out std_logic;
       MGPIO28A_OUT : out std_logic;
       MGPIO29A_OUT : out std_logic;
       MGPIO2B_OUT : out std_logic;
       MGPIO30A_OUT : out std_logic;
       MGPIO31A_OUT : out std_logic;
       MGPIO3B_OUT : out std_logic;
       MGPIO4B_OUT : out std_logic;
       MGPIO5B_OUT : out std_logic;
       MGPIO6B_OUT : out std_logic;
       MGPIO7B_OUT : out std_logic;
       MGPIO8B_OUT : out std_logic;
       MGPIO9B_OUT : out std_logic;
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT : out std_logic;
       MMUART0_DCD_MGPIO22B_OUT : out std_logic;
       MMUART0_DSR_MGPIO20B_OUT : out std_logic;
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT : out std_logic;
       MMUART0_RI_MGPIO21B_OUT : out std_logic;
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT : out std_logic;
       MMUART0_RXD_USBC_STP_MGPIO28B_OUT : out std_logic;
       MMUART0_SCK_USBC_NXT_MGPIO29B_OUT : out std_logic;
       MMUART0_TXD_USBC_DIR_MGPIO27B_OUT : out std_logic;
       MMUART1_CTS_MGPIO13B_OUT : out std_logic;
       MMUART1_DCD_MGPIO16B_OUT : out std_logic;
       MMUART1_DSR_MGPIO14B_OUT : out std_logic;
       MMUART1_DTR_MGPIO12B_OUT : out std_logic;
       MMUART1_RI_MGPIO15B_OUT : out std_logic;
       MMUART1_RTS_MGPIO11B_OUT : out std_logic;
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT : out std_logic;
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT : out std_logic;
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT : out std_logic;
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT : out std_logic;
       RGMII_MDC_RMII_MDC_OUT : out std_logic;
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT : out std_logic;
       RGMII_RX_CLK_OUT : out std_logic;
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT : out std_logic;
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT : out std_logic;
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT : out std_logic;
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT : out std_logic;
       RGMII_RXD3_USBB_DATA4_OUT : out std_logic;
       RGMII_TX_CLK_OUT : out std_logic;
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT : out std_logic;
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT : out std_logic;
       RGMII_TXD1_RMII_TXD1_USBB_STP_OUT : out std_logic;
       RGMII_TXD2_USBB_DATA5_OUT : out std_logic;
       RGMII_TXD3_USBB_DATA6_OUT : out std_logic;
       SPI0_SCK_USBA_XCLK_OUT : out std_logic;
       SPI0_SDI_USBA_DIR_MGPIO5A_OUT : out std_logic;
       SPI0_SDO_USBA_STP_MGPIO6A_OUT : out std_logic;
       SPI0_SS0_USBA_NXT_MGPIO7A_OUT : out std_logic;
       SPI0_SS1_USBA_DATA5_MGPIO8A_OUT : out std_logic;
       SPI0_SS2_USBA_DATA6_MGPIO9A_OUT : out std_logic;
       SPI0_SS3_USBA_DATA7_MGPIO10A_OUT : out std_logic;
       SPI0_SS4_MGPIO19A_OUT : out std_logic;
       SPI0_SS5_MGPIO20A_OUT : out std_logic;
       SPI0_SS6_MGPIO21A_OUT : out std_logic;
       SPI0_SS7_MGPIO22A_OUT : out std_logic;
       SPI1_SCK_OUT : out std_logic;
       SPI1_SDI_MGPIO11A_OUT : out std_logic;
       SPI1_SDO_MGPIO12A_OUT : out std_logic;
       SPI1_SS0_MGPIO13A_OUT : out std_logic;
       SPI1_SS1_MGPIO14A_OUT : out std_logic;
       SPI1_SS2_MGPIO15A_OUT : out std_logic;
       SPI1_SS3_MGPIO16A_OUT : out std_logic;
       SPI1_SS4_MGPIO17A_OUT : out std_logic;
       SPI1_SS5_MGPIO18A_OUT : out std_logic;
       SPI1_SS6_MGPIO23A_OUT : out std_logic;
       SPI1_SS7_MGPIO24A_OUT : out std_logic;
       USBC_XCLK_OUT : out std_logic;
       USBD_DATA0_OUT : out std_logic;
       USBD_DATA1_OUT : out std_logic;
       USBD_DATA2_OUT : out std_logic;
       USBD_DATA3_OUT : out std_logic;
       USBD_DATA4_OUT : out std_logic;
       USBD_DATA5_OUT : out std_logic;
       USBD_DATA6_OUT : out std_logic;
       USBD_DATA7_MGPIO23B_OUT : out std_logic;
       USBD_DIR_OUT : out std_logic;
       USBD_NXT_OUT : out std_logic;
       USBD_STP_OUT : out std_logic;
       USBD_XCLK_OUT : out std_logic;
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OE : out std_logic;
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE : out std_logic;
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OE : out std_logic;
       DM_OE : out std_logic_vector(4 downto 0);
       DRAM_DQ_OE : out std_logic_vector(35 downto 0);
       DRAM_DQS_OE : out std_logic_vector(4 downto 0);
       I2C0_SCL_USBC_DATA1_MGPIO31B_OE : out std_logic;
       I2C0_SDA_USBC_DATA0_MGPIO30B_OE : out std_logic;
       I2C1_SCL_USBA_DATA4_MGPIO1A_OE : out std_logic;
       I2C1_SDA_USBA_DATA3_MGPIO0A_OE : out std_logic;
       MGPIO0B_OE : out std_logic;
       MGPIO10B_OE : out std_logic;
       MGPIO1B_OE : out std_logic;
       MGPIO25A_OE : out std_logic;
       MGPIO26A_OE : out std_logic;
       MGPIO27A_OE : out std_logic;
       MGPIO28A_OE : out std_logic;
       MGPIO29A_OE : out std_logic;
       MGPIO2B_OE : out std_logic;
       MGPIO30A_OE : out std_logic;
       MGPIO31A_OE : out std_logic;
       MGPIO3B_OE : out std_logic;
       MGPIO4B_OE : out std_logic;
       MGPIO5B_OE : out std_logic;
       MGPIO6B_OE : out std_logic;
       MGPIO7B_OE : out std_logic;
       MGPIO8B_OE : out std_logic;
       MGPIO9B_OE : out std_logic;
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OE : out std_logic;
       MMUART0_DCD_MGPIO22B_OE : out std_logic;
       MMUART0_DSR_MGPIO20B_OE : out std_logic;
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OE : out std_logic;
       MMUART0_RI_MGPIO21B_OE : out std_logic;
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OE : out std_logic;
       MMUART0_RXD_USBC_STP_MGPIO28B_OE : out std_logic;
       MMUART0_SCK_USBC_NXT_MGPIO29B_OE : out std_logic;
       MMUART0_TXD_USBC_DIR_MGPIO27B_OE : out std_logic;
       MMUART1_CTS_MGPIO13B_OE : out std_logic;
       MMUART1_DCD_MGPIO16B_OE : out std_logic;
       MMUART1_DSR_MGPIO14B_OE : out std_logic;
       MMUART1_DTR_MGPIO12B_OE : out std_logic;
       MMUART1_RI_MGPIO15B_OE : out std_logic;
       MMUART1_RTS_MGPIO11B_OE : out std_logic;
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OE : out std_logic;
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OE : out std_logic;
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OE : out std_logic;
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE : out std_logic;
       RGMII_MDC_RMII_MDC_OE : out std_logic;
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE : out std_logic;
       RGMII_RX_CLK_OE : out std_logic;
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE : out std_logic;
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE : out std_logic;
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE : out std_logic;
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE : out std_logic;
       RGMII_RXD3_USBB_DATA4_OE : out std_logic;
       RGMII_TX_CLK_OE : out std_logic;
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE : out std_logic;
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OE : out std_logic;
       RGMII_TXD1_RMII_TXD1_USBB_STP_OE : out std_logic;
       RGMII_TXD2_USBB_DATA5_OE : out std_logic;
       RGMII_TXD3_USBB_DATA6_OE : out std_logic;
       SPI0_SCK_USBA_XCLK_OE : out std_logic;
       SPI0_SDI_USBA_DIR_MGPIO5A_OE : out std_logic;
       SPI0_SDO_USBA_STP_MGPIO6A_OE : out std_logic;
       SPI0_SS0_USBA_NXT_MGPIO7A_OE : out std_logic;
       SPI0_SS1_USBA_DATA5_MGPIO8A_OE : out std_logic;
       SPI0_SS2_USBA_DATA6_MGPIO9A_OE : out std_logic;
       SPI0_SS3_USBA_DATA7_MGPIO10A_OE : out std_logic;
       SPI0_SS4_MGPIO19A_OE : out std_logic;
       SPI0_SS5_MGPIO20A_OE : out std_logic;
       SPI0_SS6_MGPIO21A_OE : out std_logic;
       SPI0_SS7_MGPIO22A_OE : out std_logic;
       SPI1_SCK_OE : out std_logic;
       SPI1_SDI_MGPIO11A_OE : out std_logic;
       SPI1_SDO_MGPIO12A_OE : out std_logic;
       SPI1_SS0_MGPIO13A_OE : out std_logic;
       SPI1_SS1_MGPIO14A_OE : out std_logic;
       SPI1_SS2_MGPIO15A_OE : out std_logic;
       SPI1_SS3_MGPIO16A_OE : out std_logic;
       SPI1_SS4_MGPIO17A_OE : out std_logic;
       SPI1_SS5_MGPIO18A_OE : out std_logic;
       SPI1_SS6_MGPIO23A_OE : out std_logic;
       SPI1_SS7_MGPIO24A_OE : out std_logic;
       USBC_XCLK_OE : out std_logic;
       USBD_DATA0_OE : out std_logic;
       USBD_DATA1_OE : out std_logic;
       USBD_DATA2_OE : out std_logic;
       USBD_DATA3_OE : out std_logic;
       USBD_DATA4_OE : out std_logic;
       USBD_DATA5_OE : out std_logic;
       USBD_DATA6_OE : out std_logic;
       USBD_DATA7_MGPIO23B_OE : out std_logic;
       USBD_DIR_OE : out std_logic;
       USBD_NXT_OE : out std_logic;
       USBD_STP_OE : out std_logic;
       USBD_XCLK_OE : out std_logic
   );
end MSS_120;
architecture DEF_ARCH of MSS_120 is 

   attribute black_box : boolean;
   attribute black_box of DEF_ARCH : architecture is true;
   attribute ment_tsu0: string;
   attribute ment_tsu0 of DEF_ARCH : architecture is " CAN_RXBUS_F2H_SCP->CLK_BASE=1.723";
   attribute ment_tsu1: string;
   attribute ment_tsu1 of DEF_ARCH : architecture is " F2HCALIB->CLK_BASE=0.156";
   attribute ment_tsu2: string;
   attribute ment_tsu2 of DEF_ARCH : architecture is " F2H_INTERRUPT[0]->CLK_BASE=2.480";
   attribute ment_tsu3: string;
   attribute ment_tsu3 of DEF_ARCH : architecture is " F2H_INTERRUPT[10]->CLK_BASE=1.896";
   attribute ment_tsu4: string;
   attribute ment_tsu4 of DEF_ARCH : architecture is " F2H_INTERRUPT[11]->CLK_BASE=1.929";
   attribute ment_tsu5: string;
   attribute ment_tsu5 of DEF_ARCH : architecture is " F2H_INTERRUPT[12]->CLK_BASE=1.933";
   attribute ment_tsu6: string;
   attribute ment_tsu6 of DEF_ARCH : architecture is " F2H_INTERRUPT[13]->CLK_BASE=1.915";
   attribute ment_tsu7: string;
   attribute ment_tsu7 of DEF_ARCH : architecture is " F2H_INTERRUPT[14]->CLK_BASE=1.973";
   attribute ment_tsu8: string;
   attribute ment_tsu8 of DEF_ARCH : architecture is " F2H_INTERRUPT[15]->CLK_BASE=1.963";
   attribute ment_tsu9: string;
   attribute ment_tsu9 of DEF_ARCH : architecture is " F2H_INTERRUPT[1]->CLK_BASE=2.526";
   attribute ment_tsu10: string;
   attribute ment_tsu10 of DEF_ARCH : architecture is " F2H_INTERRUPT[2]->CLK_BASE=2.511";
   attribute ment_tsu11: string;
   attribute ment_tsu11 of DEF_ARCH : architecture is " F2H_INTERRUPT[3]->CLK_BASE=2.515";
   attribute ment_tsu12: string;
   attribute ment_tsu12 of DEF_ARCH : architecture is " F2H_INTERRUPT[4]->CLK_BASE=2.524";
   attribute ment_tsu13: string;
   attribute ment_tsu13 of DEF_ARCH : architecture is " F2H_INTERRUPT[5]->CLK_BASE=2.472";
   attribute ment_tsu14: string;
   attribute ment_tsu14 of DEF_ARCH : architecture is " F2H_INTERRUPT[6]->CLK_BASE=2.406";
   attribute ment_tsu15: string;
   attribute ment_tsu15 of DEF_ARCH : architecture is " F2H_INTERRUPT[7]->CLK_BASE=2.515";
   attribute ment_tsu16: string;
   attribute ment_tsu16 of DEF_ARCH : architecture is " F2H_INTERRUPT[8]->CLK_BASE=1.949";
   attribute ment_tsu17: string;
   attribute ment_tsu17 of DEF_ARCH : architecture is " F2H_INTERRUPT[9]->CLK_BASE=1.993";
   attribute ment_tsu18: string;
   attribute ment_tsu18 of DEF_ARCH : architecture is " F_FM0_ADDR[0]->CLK_BASE=0.750";
   attribute ment_tsu19: string;
   attribute ment_tsu19 of DEF_ARCH : architecture is " F_FM0_ADDR[10]->CLK_BASE=1.800";
   attribute ment_tsu20: string;
   attribute ment_tsu20 of DEF_ARCH : architecture is " F_FM0_ADDR[11]->CLK_BASE=1.886";
   attribute ment_tsu21: string;
   attribute ment_tsu21 of DEF_ARCH : architecture is " F_FM0_ADDR[12]->CLK_BASE=1.749";
   attribute ment_tsu22: string;
   attribute ment_tsu22 of DEF_ARCH : architecture is " F_FM0_ADDR[13]->CLK_BASE=1.631";
   attribute ment_tsu23: string;
   attribute ment_tsu23 of DEF_ARCH : architecture is " F_FM0_ADDR[14]->CLK_BASE=1.761";
   attribute ment_tsu24: string;
   attribute ment_tsu24 of DEF_ARCH : architecture is " F_FM0_ADDR[15]->CLK_BASE=1.763";
   attribute ment_tsu25: string;
   attribute ment_tsu25 of DEF_ARCH : architecture is " F_FM0_ADDR[16]->CLK_BASE=1.715";
   attribute ment_tsu26: string;
   attribute ment_tsu26 of DEF_ARCH : architecture is " F_FM0_ADDR[17]->CLK_BASE=1.693";
   attribute ment_tsu27: string;
   attribute ment_tsu27 of DEF_ARCH : architecture is " F_FM0_ADDR[18]->CLK_BASE=1.692";
   attribute ment_tsu28: string;
   attribute ment_tsu28 of DEF_ARCH : architecture is " F_FM0_ADDR[19]->CLK_BASE=1.453";
   attribute ment_tsu29: string;
   attribute ment_tsu29 of DEF_ARCH : architecture is " F_FM0_ADDR[1]->CLK_BASE=0.719";
   attribute ment_tsu30: string;
   attribute ment_tsu30 of DEF_ARCH : architecture is " F_FM0_ADDR[20]->CLK_BASE=1.428";
   attribute ment_tsu31: string;
   attribute ment_tsu31 of DEF_ARCH : architecture is " F_FM0_ADDR[21]->CLK_BASE=1.516";
   attribute ment_tsu32: string;
   attribute ment_tsu32 of DEF_ARCH : architecture is " F_FM0_ADDR[22]->CLK_BASE=1.742";
   attribute ment_tsu33: string;
   attribute ment_tsu33 of DEF_ARCH : architecture is " F_FM0_ADDR[23]->CLK_BASE=1.733";
   attribute ment_tsu34: string;
   attribute ment_tsu34 of DEF_ARCH : architecture is " F_FM0_ADDR[24]->CLK_BASE=1.435";
   attribute ment_tsu35: string;
   attribute ment_tsu35 of DEF_ARCH : architecture is " F_FM0_ADDR[25]->CLK_BASE=1.416";
   attribute ment_tsu36: string;
   attribute ment_tsu36 of DEF_ARCH : architecture is " F_FM0_ADDR[26]->CLK_BASE=1.460";
   attribute ment_tsu37: string;
   attribute ment_tsu37 of DEF_ARCH : architecture is " F_FM0_ADDR[27]->CLK_BASE=1.500";
   attribute ment_tsu38: string;
   attribute ment_tsu38 of DEF_ARCH : architecture is " F_FM0_ADDR[28]->CLK_BASE=1.460";
   attribute ment_tsu39: string;
   attribute ment_tsu39 of DEF_ARCH : architecture is " F_FM0_ADDR[29]->CLK_BASE=1.483";
   attribute ment_tsu40: string;
   attribute ment_tsu40 of DEF_ARCH : architecture is " F_FM0_ADDR[2]->CLK_BASE=0.493";
   attribute ment_tsu41: string;
   attribute ment_tsu41 of DEF_ARCH : architecture is " F_FM0_ADDR[30]->CLK_BASE=1.653";
   attribute ment_tsu42: string;
   attribute ment_tsu42 of DEF_ARCH : architecture is " F_FM0_ADDR[31]->CLK_BASE=1.473";
   attribute ment_tsu43: string;
   attribute ment_tsu43 of DEF_ARCH : architecture is " F_FM0_ADDR[3]->CLK_BASE=1.799";
   attribute ment_tsu44: string;
   attribute ment_tsu44 of DEF_ARCH : architecture is " F_FM0_ADDR[4]->CLK_BASE=1.706";
   attribute ment_tsu45: string;
   attribute ment_tsu45 of DEF_ARCH : architecture is " F_FM0_ADDR[5]->CLK_BASE=1.699";
   attribute ment_tsu46: string;
   attribute ment_tsu46 of DEF_ARCH : architecture is " F_FM0_ADDR[6]->CLK_BASE=1.689";
   attribute ment_tsu47: string;
   attribute ment_tsu47 of DEF_ARCH : architecture is " F_FM0_ADDR[7]->CLK_BASE=1.663";
   attribute ment_tsu48: string;
   attribute ment_tsu48 of DEF_ARCH : architecture is " F_FM0_ADDR[8]->CLK_BASE=1.728";
   attribute ment_tsu49: string;
   attribute ment_tsu49 of DEF_ARCH : architecture is " F_FM0_ADDR[9]->CLK_BASE=1.842";
   attribute ment_tsu50: string;
   attribute ment_tsu50 of DEF_ARCH : architecture is " F_FM0_MASTLOCK->CLK_BASE=0.252";
   attribute ment_tsu51: string;
   attribute ment_tsu51 of DEF_ARCH : architecture is " F_FM0_READY->CLK_BASE=0.733";
   attribute ment_tsu52: string;
   attribute ment_tsu52 of DEF_ARCH : architecture is " F_FM0_SEL->CLK_BASE=0.802";
   attribute ment_tsu53: string;
   attribute ment_tsu53 of DEF_ARCH : architecture is " F_FM0_SIZE[0]->CLK_BASE=0.632";
   attribute ment_tsu54: string;
   attribute ment_tsu54 of DEF_ARCH : architecture is " F_FM0_SIZE[1]->CLK_BASE=0.582";
   attribute ment_tsu55: string;
   attribute ment_tsu55 of DEF_ARCH : architecture is " F_FM0_TRANS1->CLK_BASE=0.839";
   attribute ment_tsu56: string;
   attribute ment_tsu56 of DEF_ARCH : architecture is " F_FM0_WDATA[0]->CLK_BASE=0.637";
   attribute ment_tsu57: string;
   attribute ment_tsu57 of DEF_ARCH : architecture is " F_FM0_WDATA[10]->CLK_BASE=0.712";
   attribute ment_tsu58: string;
   attribute ment_tsu58 of DEF_ARCH : architecture is " F_FM0_WDATA[11]->CLK_BASE=0.685";
   attribute ment_tsu59: string;
   attribute ment_tsu59 of DEF_ARCH : architecture is " F_FM0_WDATA[12]->CLK_BASE=0.705";
   attribute ment_tsu60: string;
   attribute ment_tsu60 of DEF_ARCH : architecture is " F_FM0_WDATA[13]->CLK_BASE=0.680";
   attribute ment_tsu61: string;
   attribute ment_tsu61 of DEF_ARCH : architecture is " F_FM0_WDATA[14]->CLK_BASE=0.670";
   attribute ment_tsu62: string;
   attribute ment_tsu62 of DEF_ARCH : architecture is " F_FM0_WDATA[15]->CLK_BASE=0.422";
   attribute ment_tsu63: string;
   attribute ment_tsu63 of DEF_ARCH : architecture is " F_FM0_WDATA[16]->CLK_BASE=0.574";
   attribute ment_tsu64: string;
   attribute ment_tsu64 of DEF_ARCH : architecture is " F_FM0_WDATA[17]->CLK_BASE=0.574";
   attribute ment_tsu65: string;
   attribute ment_tsu65 of DEF_ARCH : architecture is " F_FM0_WDATA[18]->CLK_BASE=0.523";
   attribute ment_tsu66: string;
   attribute ment_tsu66 of DEF_ARCH : architecture is " F_FM0_WDATA[19]->CLK_BASE=0.553";
   attribute ment_tsu67: string;
   attribute ment_tsu67 of DEF_ARCH : architecture is " F_FM0_WDATA[1]->CLK_BASE=0.653";
   attribute ment_tsu68: string;
   attribute ment_tsu68 of DEF_ARCH : architecture is " F_FM0_WDATA[20]->CLK_BASE=0.502";
   attribute ment_tsu69: string;
   attribute ment_tsu69 of DEF_ARCH : architecture is " F_FM0_WDATA[21]->CLK_BASE=0.536";
   attribute ment_tsu70: string;
   attribute ment_tsu70 of DEF_ARCH : architecture is " F_FM0_WDATA[22]->CLK_BASE=0.541";
   attribute ment_tsu71: string;
   attribute ment_tsu71 of DEF_ARCH : architecture is " F_FM0_WDATA[23]->CLK_BASE=0.554";
   attribute ment_tsu72: string;
   attribute ment_tsu72 of DEF_ARCH : architecture is " F_FM0_WDATA[24]->CLK_BASE=0.525";
   attribute ment_tsu73: string;
   attribute ment_tsu73 of DEF_ARCH : architecture is " F_FM0_WDATA[25]->CLK_BASE=0.564";
   attribute ment_tsu74: string;
   attribute ment_tsu74 of DEF_ARCH : architecture is " F_FM0_WDATA[26]->CLK_BASE=0.264";
   attribute ment_tsu75: string;
   attribute ment_tsu75 of DEF_ARCH : architecture is " F_FM0_WDATA[27]->CLK_BASE=0.550";
   attribute ment_tsu76: string;
   attribute ment_tsu76 of DEF_ARCH : architecture is " F_FM0_WDATA[28]->CLK_BASE=0.549";
   attribute ment_tsu77: string;
   attribute ment_tsu77 of DEF_ARCH : architecture is " F_FM0_WDATA[29]->CLK_BASE=0.530";
   attribute ment_tsu78: string;
   attribute ment_tsu78 of DEF_ARCH : architecture is " F_FM0_WDATA[2]->CLK_BASE=0.638";
   attribute ment_tsu79: string;
   attribute ment_tsu79 of DEF_ARCH : architecture is " F_FM0_WDATA[30]->CLK_BASE=0.533";
   attribute ment_tsu80: string;
   attribute ment_tsu80 of DEF_ARCH : architecture is " F_FM0_WDATA[31]->CLK_BASE=0.574";
   attribute ment_tsu81: string;
   attribute ment_tsu81 of DEF_ARCH : architecture is " F_FM0_WDATA[3]->CLK_BASE=0.643";
   attribute ment_tsu82: string;
   attribute ment_tsu82 of DEF_ARCH : architecture is " F_FM0_WDATA[4]->CLK_BASE=0.630";
   attribute ment_tsu83: string;
   attribute ment_tsu83 of DEF_ARCH : architecture is " F_FM0_WDATA[5]->CLK_BASE=0.691";
   attribute ment_tsu84: string;
   attribute ment_tsu84 of DEF_ARCH : architecture is " F_FM0_WDATA[6]->CLK_BASE=0.676";
   attribute ment_tsu85: string;
   attribute ment_tsu85 of DEF_ARCH : architecture is " F_FM0_WDATA[7]->CLK_BASE=0.682";
   attribute ment_tsu86: string;
   attribute ment_tsu86 of DEF_ARCH : architecture is " F_FM0_WDATA[8]->CLK_BASE=0.651";
   attribute ment_tsu87: string;
   attribute ment_tsu87 of DEF_ARCH : architecture is " F_FM0_WDATA[9]->CLK_BASE=0.692";
   attribute ment_tsu88: string;
   attribute ment_tsu88 of DEF_ARCH : architecture is " F_FM0_WRITE->CLK_BASE=0.647";
   attribute ment_tsu89: string;
   attribute ment_tsu89 of DEF_ARCH : architecture is " F_FM1_ADDR[0]->CLK_BASE=0.460";
   attribute ment_tsu90: string;
   attribute ment_tsu90 of DEF_ARCH : architecture is " F_FM1_ADDR[10]->CLK_BASE=1.118";
   attribute ment_tsu91: string;
   attribute ment_tsu91 of DEF_ARCH : architecture is " F_FM1_ADDR[11]->CLK_BASE=1.087";
   attribute ment_tsu92: string;
   attribute ment_tsu92 of DEF_ARCH : architecture is " F_FM1_ADDR[12]->CLK_BASE=1.052";
   attribute ment_tsu93: string;
   attribute ment_tsu93 of DEF_ARCH : architecture is " F_FM1_ADDR[13]->CLK_BASE=1.219";
   attribute ment_tsu94: string;
   attribute ment_tsu94 of DEF_ARCH : architecture is " F_FM1_ADDR[14]->CLK_BASE=1.117";
   attribute ment_tsu95: string;
   attribute ment_tsu95 of DEF_ARCH : architecture is " F_FM1_ADDR[15]->CLK_BASE=1.029";
   attribute ment_tsu96: string;
   attribute ment_tsu96 of DEF_ARCH : architecture is " F_FM1_ADDR[16]->CLK_BASE=1.074";
   attribute ment_tsu97: string;
   attribute ment_tsu97 of DEF_ARCH : architecture is " F_FM1_ADDR[17]->CLK_BASE=1.091";
   attribute ment_tsu98: string;
   attribute ment_tsu98 of DEF_ARCH : architecture is " F_FM1_ADDR[18]->CLK_BASE=1.041";
   attribute ment_tsu99: string;
   attribute ment_tsu99 of DEF_ARCH : architecture is " F_FM1_ADDR[19]->CLK_BASE=1.156";
   attribute ment_tsu100: string;
   attribute ment_tsu100 of DEF_ARCH : architecture is " F_FM1_ADDR[1]->CLK_BASE=0.452";
   attribute ment_tsu101: string;
   attribute ment_tsu101 of DEF_ARCH : architecture is " F_FM1_ADDR[20]->CLK_BASE=1.031";
   attribute ment_tsu102: string;
   attribute ment_tsu102 of DEF_ARCH : architecture is " F_FM1_ADDR[21]->CLK_BASE=0.897";
   attribute ment_tsu103: string;
   attribute ment_tsu103 of DEF_ARCH : architecture is " F_FM1_ADDR[22]->CLK_BASE=0.858";
   attribute ment_tsu104: string;
   attribute ment_tsu104 of DEF_ARCH : architecture is " F_FM1_ADDR[23]->CLK_BASE=1.058";
   attribute ment_tsu105: string;
   attribute ment_tsu105 of DEF_ARCH : architecture is " F_FM1_ADDR[24]->CLK_BASE=1.103";
   attribute ment_tsu106: string;
   attribute ment_tsu106 of DEF_ARCH : architecture is " F_FM1_ADDR[25]->CLK_BASE=0.891";
   attribute ment_tsu107: string;
   attribute ment_tsu107 of DEF_ARCH : architecture is " F_FM1_ADDR[26]->CLK_BASE=0.905";
   attribute ment_tsu108: string;
   attribute ment_tsu108 of DEF_ARCH : architecture is " F_FM1_ADDR[27]->CLK_BASE=0.941";
   attribute ment_tsu109: string;
   attribute ment_tsu109 of DEF_ARCH : architecture is " F_FM1_ADDR[28]->CLK_BASE=0.812";
   attribute ment_tsu110: string;
   attribute ment_tsu110 of DEF_ARCH : architecture is " F_FM1_ADDR[29]->CLK_BASE=0.794";
   attribute ment_tsu111: string;
   attribute ment_tsu111 of DEF_ARCH : architecture is " F_FM1_ADDR[2]->CLK_BASE=0.304";
   attribute ment_tsu112: string;
   attribute ment_tsu112 of DEF_ARCH : architecture is " F_FM1_ADDR[30]->CLK_BASE=1.001";
   attribute ment_tsu113: string;
   attribute ment_tsu113 of DEF_ARCH : architecture is " F_FM1_ADDR[31]->CLK_BASE=0.826";
   attribute ment_tsu114: string;
   attribute ment_tsu114 of DEF_ARCH : architecture is " F_FM1_ADDR[3]->CLK_BASE=1.146";
   attribute ment_tsu115: string;
   attribute ment_tsu115 of DEF_ARCH : architecture is " F_FM1_ADDR[4]->CLK_BASE=1.157";
   attribute ment_tsu116: string;
   attribute ment_tsu116 of DEF_ARCH : architecture is " F_FM1_ADDR[5]->CLK_BASE=1.460";
   attribute ment_tsu117: string;
   attribute ment_tsu117 of DEF_ARCH : architecture is " F_FM1_ADDR[6]->CLK_BASE=1.428";
   attribute ment_tsu118: string;
   attribute ment_tsu118 of DEF_ARCH : architecture is " F_FM1_ADDR[7]->CLK_BASE=1.140";
   attribute ment_tsu119: string;
   attribute ment_tsu119 of DEF_ARCH : architecture is " F_FM1_ADDR[8]->CLK_BASE=1.152";
   attribute ment_tsu120: string;
   attribute ment_tsu120 of DEF_ARCH : architecture is " F_FM1_ADDR[9]->CLK_BASE=1.114";
   attribute ment_tsu121: string;
   attribute ment_tsu121 of DEF_ARCH : architecture is " F_FM1_ENABLE->CLK_BASE=0.871";
   attribute ment_tsu122: string;
   attribute ment_tsu122 of DEF_ARCH : architecture is " F_FM1_SEL->CLK_BASE=0.757";
   attribute ment_tsu123: string;
   attribute ment_tsu123 of DEF_ARCH : architecture is " F_FM1_WDATA[0]->CLK_BASE=0.629";
   attribute ment_tsu124: string;
   attribute ment_tsu124 of DEF_ARCH : architecture is " F_FM1_WDATA[10]->CLK_BASE=0.755";
   attribute ment_tsu125: string;
   attribute ment_tsu125 of DEF_ARCH : architecture is " F_FM1_WDATA[11]->CLK_BASE=0.633";
   attribute ment_tsu126: string;
   attribute ment_tsu126 of DEF_ARCH : architecture is " F_FM1_WDATA[12]->CLK_BASE=0.691";
   attribute ment_tsu127: string;
   attribute ment_tsu127 of DEF_ARCH : architecture is " F_FM1_WDATA[13]->CLK_BASE=0.403";
   attribute ment_tsu128: string;
   attribute ment_tsu128 of DEF_ARCH : architecture is " F_FM1_WDATA[14]->CLK_BASE=0.705";
   attribute ment_tsu129: string;
   attribute ment_tsu129 of DEF_ARCH : architecture is " F_FM1_WDATA[15]->CLK_BASE=0.561";
   attribute ment_tsu130: string;
   attribute ment_tsu130 of DEF_ARCH : architecture is " F_FM1_WDATA[16]->CLK_BASE=0.616";
   attribute ment_tsu131: string;
   attribute ment_tsu131 of DEF_ARCH : architecture is " F_FM1_WDATA[17]->CLK_BASE=0.724";
   attribute ment_tsu132: string;
   attribute ment_tsu132 of DEF_ARCH : architecture is " F_FM1_WDATA[18]->CLK_BASE=0.606";
   attribute ment_tsu133: string;
   attribute ment_tsu133 of DEF_ARCH : architecture is " F_FM1_WDATA[19]->CLK_BASE=0.662";
   attribute ment_tsu134: string;
   attribute ment_tsu134 of DEF_ARCH : architecture is " F_FM1_WDATA[1]->CLK_BASE=0.687";
   attribute ment_tsu135: string;
   attribute ment_tsu135 of DEF_ARCH : architecture is " F_FM1_WDATA[20]->CLK_BASE=0.278";
   attribute ment_tsu136: string;
   attribute ment_tsu136 of DEF_ARCH : architecture is " F_FM1_WDATA[21]->CLK_BASE=0.619";
   attribute ment_tsu137: string;
   attribute ment_tsu137 of DEF_ARCH : architecture is " F_FM1_WDATA[22]->CLK_BASE=0.566";
   attribute ment_tsu138: string;
   attribute ment_tsu138 of DEF_ARCH : architecture is " F_FM1_WDATA[23]->CLK_BASE=0.302";
   attribute ment_tsu139: string;
   attribute ment_tsu139 of DEF_ARCH : architecture is " F_FM1_WDATA[24]->CLK_BASE=0.535";
   attribute ment_tsu140: string;
   attribute ment_tsu140 of DEF_ARCH : architecture is " F_FM1_WDATA[25]->CLK_BASE=0.689";
   attribute ment_tsu141: string;
   attribute ment_tsu141 of DEF_ARCH : architecture is " F_FM1_WDATA[26]->CLK_BASE=0.645";
   attribute ment_tsu142: string;
   attribute ment_tsu142 of DEF_ARCH : architecture is " F_FM1_WDATA[27]->CLK_BASE=0.584";
   attribute ment_tsu143: string;
   attribute ment_tsu143 of DEF_ARCH : architecture is " F_FM1_WDATA[28]->CLK_BASE=0.697";
   attribute ment_tsu144: string;
   attribute ment_tsu144 of DEF_ARCH : architecture is " F_FM1_WDATA[29]->CLK_BASE=0.655";
   attribute ment_tsu145: string;
   attribute ment_tsu145 of DEF_ARCH : architecture is " F_FM1_WDATA[2]->CLK_BASE=0.708";
   attribute ment_tsu146: string;
   attribute ment_tsu146 of DEF_ARCH : architecture is " F_FM1_WDATA[30]->CLK_BASE=0.669";
   attribute ment_tsu147: string;
   attribute ment_tsu147 of DEF_ARCH : architecture is " F_FM1_WDATA[31]->CLK_BASE=0.613";
   attribute ment_tsu148: string;
   attribute ment_tsu148 of DEF_ARCH : architecture is " F_FM1_WDATA[3]->CLK_BASE=0.627";
   attribute ment_tsu149: string;
   attribute ment_tsu149 of DEF_ARCH : architecture is " F_FM1_WDATA[4]->CLK_BASE=0.648";
   attribute ment_tsu150: string;
   attribute ment_tsu150 of DEF_ARCH : architecture is " F_FM1_WDATA[5]->CLK_BASE=0.288";
   attribute ment_tsu151: string;
   attribute ment_tsu151 of DEF_ARCH : architecture is " F_FM1_WDATA[6]->CLK_BASE=0.671";
   attribute ment_tsu152: string;
   attribute ment_tsu152 of DEF_ARCH : architecture is " F_FM1_WDATA[7]->CLK_BASE=0.650";
   attribute ment_tsu153: string;
   attribute ment_tsu153 of DEF_ARCH : architecture is " F_FM1_WDATA[8]->CLK_BASE=0.627";
   attribute ment_tsu154: string;
   attribute ment_tsu154 of DEF_ARCH : architecture is " F_FM1_WDATA[9]->CLK_BASE=0.354";
   attribute ment_tsu155: string;
   attribute ment_tsu155 of DEF_ARCH : architecture is " F_FM1_WRITE->CLK_BASE=0.784";
   attribute ment_tsu156: string;
   attribute ment_tsu156 of DEF_ARCH : architecture is " F_HM0_RDATA[0]->CLK_BASE=0.550";
   attribute ment_tsu157: string;
   attribute ment_tsu157 of DEF_ARCH : architecture is " F_HM0_RDATA[10]->CLK_BASE=0.564";
   attribute ment_tsu158: string;
   attribute ment_tsu158 of DEF_ARCH : architecture is " F_HM0_RDATA[11]->CLK_BASE=0.524";
   attribute ment_tsu159: string;
   attribute ment_tsu159 of DEF_ARCH : architecture is " F_HM0_RDATA[12]->CLK_BASE=0.512";
   attribute ment_tsu160: string;
   attribute ment_tsu160 of DEF_ARCH : architecture is " F_HM0_RDATA[13]->CLK_BASE=0.525";
   attribute ment_tsu161: string;
   attribute ment_tsu161 of DEF_ARCH : architecture is " F_HM0_RDATA[14]->CLK_BASE=0.516";
   attribute ment_tsu162: string;
   attribute ment_tsu162 of DEF_ARCH : architecture is " F_HM0_RDATA[15]->CLK_BASE=0.539";
   attribute ment_tsu163: string;
   attribute ment_tsu163 of DEF_ARCH : architecture is " F_HM0_RDATA[16]->CLK_BASE=0.487";
   attribute ment_tsu164: string;
   attribute ment_tsu164 of DEF_ARCH : architecture is " F_HM0_RDATA[17]->CLK_BASE=0.494";
   attribute ment_tsu165: string;
   attribute ment_tsu165 of DEF_ARCH : architecture is " F_HM0_RDATA[18]->CLK_BASE=0.521";
   attribute ment_tsu166: string;
   attribute ment_tsu166 of DEF_ARCH : architecture is " F_HM0_RDATA[19]->CLK_BASE=0.553";
   attribute ment_tsu167: string;
   attribute ment_tsu167 of DEF_ARCH : architecture is " F_HM0_RDATA[1]->CLK_BASE=0.596";
   attribute ment_tsu168: string;
   attribute ment_tsu168 of DEF_ARCH : architecture is " F_HM0_RDATA[20]->CLK_BASE=0.516";
   attribute ment_tsu169: string;
   attribute ment_tsu169 of DEF_ARCH : architecture is " F_HM0_RDATA[21]->CLK_BASE=0.526";
   attribute ment_tsu170: string;
   attribute ment_tsu170 of DEF_ARCH : architecture is " F_HM0_RDATA[22]->CLK_BASE=0.513";
   attribute ment_tsu171: string;
   attribute ment_tsu171 of DEF_ARCH : architecture is " F_HM0_RDATA[23]->CLK_BASE=0.537";
   attribute ment_tsu172: string;
   attribute ment_tsu172 of DEF_ARCH : architecture is " F_HM0_RDATA[24]->CLK_BASE=0.460";
   attribute ment_tsu173: string;
   attribute ment_tsu173 of DEF_ARCH : architecture is " F_HM0_RDATA[25]->CLK_BASE=0.574";
   attribute ment_tsu174: string;
   attribute ment_tsu174 of DEF_ARCH : architecture is " F_HM0_RDATA[26]->CLK_BASE=0.508";
   attribute ment_tsu175: string;
   attribute ment_tsu175 of DEF_ARCH : architecture is " F_HM0_RDATA[27]->CLK_BASE=0.521";
   attribute ment_tsu176: string;
   attribute ment_tsu176 of DEF_ARCH : architecture is " F_HM0_RDATA[28]->CLK_BASE=0.495";
   attribute ment_tsu177: string;
   attribute ment_tsu177 of DEF_ARCH : architecture is " F_HM0_RDATA[29]->CLK_BASE=0.500";
   attribute ment_tsu178: string;
   attribute ment_tsu178 of DEF_ARCH : architecture is " F_HM0_RDATA[2]->CLK_BASE=0.576";
   attribute ment_tsu179: string;
   attribute ment_tsu179 of DEF_ARCH : architecture is " F_HM0_RDATA[30]->CLK_BASE=0.516";
   attribute ment_tsu180: string;
   attribute ment_tsu180 of DEF_ARCH : architecture is " F_HM0_RDATA[31]->CLK_BASE=0.466";
   attribute ment_tsu181: string;
   attribute ment_tsu181 of DEF_ARCH : architecture is " F_HM0_RDATA[3]->CLK_BASE=0.598";
   attribute ment_tsu182: string;
   attribute ment_tsu182 of DEF_ARCH : architecture is " F_HM0_RDATA[4]->CLK_BASE=0.554";
   attribute ment_tsu183: string;
   attribute ment_tsu183 of DEF_ARCH : architecture is " F_HM0_RDATA[5]->CLK_BASE=0.580";
   attribute ment_tsu184: string;
   attribute ment_tsu184 of DEF_ARCH : architecture is " F_HM0_RDATA[6]->CLK_BASE=0.556";
   attribute ment_tsu185: string;
   attribute ment_tsu185 of DEF_ARCH : architecture is " F_HM0_RDATA[7]->CLK_BASE=0.589";
   attribute ment_tsu186: string;
   attribute ment_tsu186 of DEF_ARCH : architecture is " F_HM0_RDATA[8]->CLK_BASE=0.548";
   attribute ment_tsu187: string;
   attribute ment_tsu187 of DEF_ARCH : architecture is " F_HM0_RDATA[9]->CLK_BASE=0.533";
   attribute ment_tsu188: string;
   attribute ment_tsu188 of DEF_ARCH : architecture is " F_HM0_READY->CLK_BASE=0.779";
   attribute ment_tsu189: string;
   attribute ment_tsu189 of DEF_ARCH : architecture is " F_HM0_RESP->CLK_BASE=0.764";
   attribute ment_tsu190: string;
   attribute ment_tsu190 of DEF_ARCH : architecture is " F_HM1_RDATA[0]->CLK_BASE=0.489";
   attribute ment_tsu191: string;
   attribute ment_tsu191 of DEF_ARCH : architecture is " F_HM1_RDATA[10]->CLK_BASE=0.542";
   attribute ment_tsu192: string;
   attribute ment_tsu192 of DEF_ARCH : architecture is " F_HM1_RDATA[11]->CLK_BASE=0.533";
   attribute ment_tsu193: string;
   attribute ment_tsu193 of DEF_ARCH : architecture is " F_HM1_RDATA[12]->CLK_BASE=0.559";
   attribute ment_tsu194: string;
   attribute ment_tsu194 of DEF_ARCH : architecture is " F_HM1_RDATA[13]->CLK_BASE=0.521";
   attribute ment_tsu195: string;
   attribute ment_tsu195 of DEF_ARCH : architecture is " F_HM1_RDATA[14]->CLK_BASE=0.542";
   attribute ment_tsu196: string;
   attribute ment_tsu196 of DEF_ARCH : architecture is " F_HM1_RDATA[15]->CLK_BASE=0.539";
   attribute ment_tsu197: string;
   attribute ment_tsu197 of DEF_ARCH : architecture is " F_HM1_RDATA[16]->CLK_BASE=0.548";
   attribute ment_tsu198: string;
   attribute ment_tsu198 of DEF_ARCH : architecture is " F_HM1_RDATA[17]->CLK_BASE=0.531";
   attribute ment_tsu199: string;
   attribute ment_tsu199 of DEF_ARCH : architecture is " F_HM1_RDATA[18]->CLK_BASE=0.498";
   attribute ment_tsu200: string;
   attribute ment_tsu200 of DEF_ARCH : architecture is " F_HM1_RDATA[19]->CLK_BASE=0.503";
   attribute ment_tsu201: string;
   attribute ment_tsu201 of DEF_ARCH : architecture is " F_HM1_RDATA[1]->CLK_BASE=0.517";
   attribute ment_tsu202: string;
   attribute ment_tsu202 of DEF_ARCH : architecture is " F_HM1_RDATA[20]->CLK_BASE=0.516";
   attribute ment_tsu203: string;
   attribute ment_tsu203 of DEF_ARCH : architecture is " F_HM1_RDATA[21]->CLK_BASE=0.489";
   attribute ment_tsu204: string;
   attribute ment_tsu204 of DEF_ARCH : architecture is " F_HM1_RDATA[22]->CLK_BASE=0.506";
   attribute ment_tsu205: string;
   attribute ment_tsu205 of DEF_ARCH : architecture is " F_HM1_RDATA[23]->CLK_BASE=0.510";
   attribute ment_tsu206: string;
   attribute ment_tsu206 of DEF_ARCH : architecture is " F_HM1_RDATA[24]->CLK_BASE=0.519";
   attribute ment_tsu207: string;
   attribute ment_tsu207 of DEF_ARCH : architecture is " F_HM1_RDATA[25]->CLK_BASE=0.508";
   attribute ment_tsu208: string;
   attribute ment_tsu208 of DEF_ARCH : architecture is " F_HM1_RDATA[26]->CLK_BASE=0.539";
   attribute ment_tsu209: string;
   attribute ment_tsu209 of DEF_ARCH : architecture is " F_HM1_RDATA[27]->CLK_BASE=0.525";
   attribute ment_tsu210: string;
   attribute ment_tsu210 of DEF_ARCH : architecture is " F_HM1_RDATA[28]->CLK_BASE=0.509";
   attribute ment_tsu211: string;
   attribute ment_tsu211 of DEF_ARCH : architecture is " F_HM1_RDATA[29]->CLK_BASE=0.520";
   attribute ment_tsu212: string;
   attribute ment_tsu212 of DEF_ARCH : architecture is " F_HM1_RDATA[2]->CLK_BASE=0.523";
   attribute ment_tsu213: string;
   attribute ment_tsu213 of DEF_ARCH : architecture is " F_HM1_RDATA[30]->CLK_BASE=0.547";
   attribute ment_tsu214: string;
   attribute ment_tsu214 of DEF_ARCH : architecture is " F_HM1_RDATA[31]->CLK_BASE=0.526";
   attribute ment_tsu215: string;
   attribute ment_tsu215 of DEF_ARCH : architecture is " F_HM1_RDATA[3]->CLK_BASE=0.533";
   attribute ment_tsu216: string;
   attribute ment_tsu216 of DEF_ARCH : architecture is " F_HM1_RDATA[4]->CLK_BASE=0.502";
   attribute ment_tsu217: string;
   attribute ment_tsu217 of DEF_ARCH : architecture is " F_HM1_RDATA[5]->CLK_BASE=0.505";
   attribute ment_tsu218: string;
   attribute ment_tsu218 of DEF_ARCH : architecture is " F_HM1_RDATA[6]->CLK_BASE=0.508";
   attribute ment_tsu219: string;
   attribute ment_tsu219 of DEF_ARCH : architecture is " F_HM1_RDATA[7]->CLK_BASE=0.497";
   attribute ment_tsu220: string;
   attribute ment_tsu220 of DEF_ARCH : architecture is " F_HM1_RDATA[8]->CLK_BASE=0.561";
   attribute ment_tsu221: string;
   attribute ment_tsu221 of DEF_ARCH : architecture is " F_HM1_RDATA[9]->CLK_BASE=0.522";
   attribute ment_tsu222: string;
   attribute ment_tsu222 of DEF_ARCH : architecture is " F_HM1_READY->CLK_BASE=0.831";
   attribute ment_tsu223: string;
   attribute ment_tsu223 of DEF_ARCH : architecture is " F_HM1_RESP->CLK_BASE=0.816";
   attribute ment_tsu224: string;
   attribute ment_tsu224 of DEF_ARCH : architecture is " I2C0_SDA_F2H_SCP->I2C0_SCL_F2H_SCP=0.024";
   attribute ment_tsu225: string;
   attribute ment_tsu225 of DEF_ARCH : architecture is " I2C1_SDA_F2H_SCP->I2C1_SCL_F2H_SCP=-0.023";
   attribute ment_tsu226: string;
   attribute ment_tsu226 of DEF_ARCH : architecture is " MDDR_FABRIC_PADDR[10]->CLK_MDDR_APB=0.413";
   attribute ment_tsu227: string;
   attribute ment_tsu227 of DEF_ARCH : architecture is " MDDR_FABRIC_PADDR[2]->CLK_MDDR_APB=0.392";
   attribute ment_tsu228: string;
   attribute ment_tsu228 of DEF_ARCH : architecture is " MDDR_FABRIC_PADDR[3]->CLK_MDDR_APB=0.343";
   attribute ment_tsu229: string;
   attribute ment_tsu229 of DEF_ARCH : architecture is " MDDR_FABRIC_PADDR[4]->CLK_MDDR_APB=0.410";
   attribute ment_tsu230: string;
   attribute ment_tsu230 of DEF_ARCH : architecture is " MDDR_FABRIC_PADDR[5]->CLK_MDDR_APB=0.181";
   attribute ment_tsu231: string;
   attribute ment_tsu231 of DEF_ARCH : architecture is " MDDR_FABRIC_PADDR[6]->CLK_MDDR_APB=0.257";
   attribute ment_tsu232: string;
   attribute ment_tsu232 of DEF_ARCH : architecture is " MDDR_FABRIC_PADDR[7]->CLK_MDDR_APB=0.186";
   attribute ment_tsu233: string;
   attribute ment_tsu233 of DEF_ARCH : architecture is " MDDR_FABRIC_PADDR[8]->CLK_MDDR_APB=0.312";
   attribute ment_tsu234: string;
   attribute ment_tsu234 of DEF_ARCH : architecture is " MDDR_FABRIC_PADDR[9]->CLK_MDDR_APB=0.364";
   attribute ment_tsu235: string;
   attribute ment_tsu235 of DEF_ARCH : architecture is " MDDR_FABRIC_PENABLE->CLK_MDDR_APB=0.332";
   attribute ment_tsu236: string;
   attribute ment_tsu236 of DEF_ARCH : architecture is " MDDR_FABRIC_PSEL->CLK_MDDR_APB=0.396";
   attribute ment_tsu237: string;
   attribute ment_tsu237 of DEF_ARCH : architecture is " MDDR_FABRIC_PWDATA[0]->CLK_MDDR_APB=0.408";
   attribute ment_tsu238: string;
   attribute ment_tsu238 of DEF_ARCH : architecture is " MDDR_FABRIC_PWDATA[10]->CLK_MDDR_APB=-0.218";
   attribute ment_tsu239: string;
   attribute ment_tsu239 of DEF_ARCH : architecture is " MDDR_FABRIC_PWDATA[11]->CLK_MDDR_APB=-0.100";
   attribute ment_tsu240: string;
   attribute ment_tsu240 of DEF_ARCH : architecture is " MDDR_FABRIC_PWDATA[12]->CLK_MDDR_APB=-0.322";
   attribute ment_tsu241: string;
   attribute ment_tsu241 of DEF_ARCH : architecture is " MDDR_FABRIC_PWDATA[13]->CLK_MDDR_APB=-0.409";
   attribute ment_tsu242: string;
   attribute ment_tsu242 of DEF_ARCH : architecture is " MDDR_FABRIC_PWDATA[14]->CLK_MDDR_APB=-0.404";
   attribute ment_tsu243: string;
   attribute ment_tsu243 of DEF_ARCH : architecture is " MDDR_FABRIC_PWDATA[15]->CLK_MDDR_APB=-0.391";
   attribute ment_tsu244: string;
   attribute ment_tsu244 of DEF_ARCH : architecture is " MDDR_FABRIC_PWDATA[1]->CLK_MDDR_APB=0.466";
   attribute ment_tsu245: string;
   attribute ment_tsu245 of DEF_ARCH : architecture is " MDDR_FABRIC_PWDATA[2]->CLK_MDDR_APB=-0.129";
   attribute ment_tsu246: string;
   attribute ment_tsu246 of DEF_ARCH : architecture is " MDDR_FABRIC_PWDATA[3]->CLK_MDDR_APB=-0.254";
   attribute ment_tsu247: string;
   attribute ment_tsu247 of DEF_ARCH : architecture is " MDDR_FABRIC_PWDATA[4]->CLK_MDDR_APB=-0.233";
   attribute ment_tsu248: string;
   attribute ment_tsu248 of DEF_ARCH : architecture is " MDDR_FABRIC_PWDATA[5]->CLK_MDDR_APB=-0.377";
   attribute ment_tsu249: string;
   attribute ment_tsu249 of DEF_ARCH : architecture is " MDDR_FABRIC_PWDATA[6]->CLK_MDDR_APB=-0.431";
   attribute ment_tsu250: string;
   attribute ment_tsu250 of DEF_ARCH : architecture is " MDDR_FABRIC_PWDATA[7]->CLK_MDDR_APB=-0.078";
   attribute ment_tsu251: string;
   attribute ment_tsu251 of DEF_ARCH : architecture is " MDDR_FABRIC_PWDATA[8]->CLK_MDDR_APB=-0.408";
   attribute ment_tsu252: string;
   attribute ment_tsu252 of DEF_ARCH : architecture is " MDDR_FABRIC_PWDATA[9]->CLK_MDDR_APB=-0.182";
   attribute ment_tsu253: string;
   attribute ment_tsu253 of DEF_ARCH : architecture is " MDDR_FABRIC_PWRITE->CLK_MDDR_APB=0.160";
   attribute ment_tsu254: string;
   attribute ment_tsu254 of DEF_ARCH : architecture is " MGPIO0A_F2H_GPIN->CLK_BASE=1.319";
   attribute ment_tsu255: string;
   attribute ment_tsu255 of DEF_ARCH : architecture is " MGPIO10A_F2H_GPIN->CLK_BASE=1.325";
   attribute ment_tsu256: string;
   attribute ment_tsu256 of DEF_ARCH : architecture is " MGPIO11A_F2H_GPIN->CLK_BASE=1.140";
   attribute ment_tsu257: string;
   attribute ment_tsu257 of DEF_ARCH : architecture is " MGPIO11B_F2H_GPIN->CLK_BASE=1.346";
   attribute ment_tsu258: string;
   attribute ment_tsu258 of DEF_ARCH : architecture is " MGPIO12A_F2H_GPIN->CLK_BASE=1.104";
   attribute ment_tsu259: string;
   attribute ment_tsu259 of DEF_ARCH : architecture is " MGPIO13A_F2H_GPIN->CLK_BASE=1.270";
   attribute ment_tsu260: string;
   attribute ment_tsu260 of DEF_ARCH : architecture is " MGPIO14A_F2H_GPIN->CLK_BASE=1.155";
   attribute ment_tsu261: string;
   attribute ment_tsu261 of DEF_ARCH : architecture is " MGPIO15A_F2H_GPIN->CLK_BASE=0.944";
   attribute ment_tsu262: string;
   attribute ment_tsu262 of DEF_ARCH : architecture is " MGPIO16A_F2H_GPIN->CLK_BASE=1.131";
   attribute ment_tsu263: string;
   attribute ment_tsu263 of DEF_ARCH : architecture is " MGPIO17B_F2H_GPIN->CLK_BASE=0.955";
   attribute ment_tsu264: string;
   attribute ment_tsu264 of DEF_ARCH : architecture is " MGPIO18B_F2H_GPIN->CLK_BASE=1.191";
   attribute ment_tsu265: string;
   attribute ment_tsu265 of DEF_ARCH : architecture is " MGPIO19B_F2H_GPIN->CLK_BASE=1.338";
   attribute ment_tsu266: string;
   attribute ment_tsu266 of DEF_ARCH : architecture is " MGPIO1A_F2H_GPIN->CLK_BASE=1.452";
   attribute ment_tsu267: string;
   attribute ment_tsu267 of DEF_ARCH : architecture is " MGPIO20B_F2H_GPIN->CLK_BASE=1.236";
   attribute ment_tsu268: string;
   attribute ment_tsu268 of DEF_ARCH : architecture is " MGPIO21B_F2H_GPIN->CLK_BASE=1.012";
   attribute ment_tsu269: string;
   attribute ment_tsu269 of DEF_ARCH : architecture is " MGPIO22B_F2H_GPIN->CLK_BASE=1.321";
   attribute ment_tsu270: string;
   attribute ment_tsu270 of DEF_ARCH : architecture is " MGPIO24B_F2H_GPIN->CLK_BASE=1.238";
   attribute ment_tsu271: string;
   attribute ment_tsu271 of DEF_ARCH : architecture is " MGPIO25B_F2H_GPIN->CLK_BASE=1.261";
   attribute ment_tsu272: string;
   attribute ment_tsu272 of DEF_ARCH : architecture is " MGPIO26B_F2H_GPIN->CLK_BASE=1.508";
   attribute ment_tsu273: string;
   attribute ment_tsu273 of DEF_ARCH : architecture is " MGPIO27B_F2H_GPIN->CLK_BASE=1.226";
   attribute ment_tsu274: string;
   attribute ment_tsu274 of DEF_ARCH : architecture is " MGPIO28B_F2H_GPIN->CLK_BASE=1.482";
   attribute ment_tsu275: string;
   attribute ment_tsu275 of DEF_ARCH : architecture is " MGPIO29B_F2H_GPIN->CLK_BASE=1.702";
   attribute ment_tsu276: string;
   attribute ment_tsu276 of DEF_ARCH : architecture is " MGPIO2A_F2H_GPIN->CLK_BASE=1.057";
   attribute ment_tsu277: string;
   attribute ment_tsu277 of DEF_ARCH : architecture is " MGPIO30B_F2H_GPIN->CLK_BASE=1.306";
   attribute ment_tsu278: string;
   attribute ment_tsu278 of DEF_ARCH : architecture is " MGPIO31B_F2H_GPIN->CLK_BASE=1.288";
   attribute ment_tsu279: string;
   attribute ment_tsu279 of DEF_ARCH : architecture is " MGPIO3A_F2H_GPIN->CLK_BASE=1.444";
   attribute ment_tsu280: string;
   attribute ment_tsu280 of DEF_ARCH : architecture is " MGPIO4A_F2H_GPIN->CLK_BASE=1.347";
   attribute ment_tsu281: string;
   attribute ment_tsu281 of DEF_ARCH : architecture is " MGPIO5A_F2H_GPIN->CLK_BASE=1.267";
   attribute ment_tsu282: string;
   attribute ment_tsu282 of DEF_ARCH : architecture is " MGPIO6A_F2H_GPIN->CLK_BASE=1.049";
   attribute ment_tsu283: string;
   attribute ment_tsu283 of DEF_ARCH : architecture is " MGPIO7A_F2H_GPIN->CLK_BASE=1.322";
   attribute ment_tsu284: string;
   attribute ment_tsu284 of DEF_ARCH : architecture is " MGPIO8A_F2H_GPIN->CLK_BASE=1.014";
   attribute ment_tsu285: string;
   attribute ment_tsu285 of DEF_ARCH : architecture is " MGPIO9A_F2H_GPIN->CLK_BASE=1.124";
   attribute ment_tsu286: string;
   attribute ment_tsu286 of DEF_ARCH : architecture is " MMUART0_CTS_F2H_SCP->CLK_BASE=1.349";
   attribute ment_tsu287: string;
   attribute ment_tsu287 of DEF_ARCH : architecture is " MMUART0_DCD_F2H_SCP->CLK_BASE=1.114";
   attribute ment_tsu288: string;
   attribute ment_tsu288 of DEF_ARCH : architecture is " MMUART0_DSR_F2H_SCP->CLK_BASE=1.077";
   attribute ment_tsu289: string;
   attribute ment_tsu289 of DEF_ARCH : architecture is " MMUART0_RI_F2H_SCP->CLK_BASE=1.194";
   attribute ment_tsu290: string;
   attribute ment_tsu290 of DEF_ARCH : architecture is " MMUART0_RXD_F2H_SCP->CLK_BASE=0.969";
   attribute ment_tsu291: string;
   attribute ment_tsu291 of DEF_ARCH : architecture is " MMUART0_SCK_F2H_SCP->CLK_BASE=1.024";
   attribute ment_tsu292: string;
   attribute ment_tsu292 of DEF_ARCH : architecture is " MMUART0_TXD_F2H_SCP->CLK_BASE=0.955";
   attribute ment_tsu293: string;
   attribute ment_tsu293 of DEF_ARCH : architecture is " MMUART1_CTS_F2H_SCP->CLK_BASE=2.033";
   attribute ment_tsu294: string;
   attribute ment_tsu294 of DEF_ARCH : architecture is " MMUART1_DCD_F2H_SCP->CLK_BASE=2.002";
   attribute ment_tsu295: string;
   attribute ment_tsu295 of DEF_ARCH : architecture is " MMUART1_DSR_F2H_SCP->CLK_BASE=2.133";
   attribute ment_tsu296: string;
   attribute ment_tsu296 of DEF_ARCH : architecture is " MMUART1_RI_F2H_SCP->CLK_BASE=1.812";
   attribute ment_tsu297: string;
   attribute ment_tsu297 of DEF_ARCH : architecture is " MMUART1_RXD_F2H_SCP->CLK_BASE=2.178";
   attribute ment_tsu298: string;
   attribute ment_tsu298 of DEF_ARCH : architecture is " MMUART1_SCK_F2H_SCP->CLK_BASE=1.959";
   attribute ment_tsu299: string;
   attribute ment_tsu299 of DEF_ARCH : architecture is " MMUART1_TXD_F2H_SCP->CLK_BASE=1.964";
   attribute ment_tsu300: string;
   attribute ment_tsu300 of DEF_ARCH : architecture is " SMBALERT_NI0->I2C0_SCL_F2H_SCP=-0.760";
   attribute ment_tsu301: string;
   attribute ment_tsu301 of DEF_ARCH : architecture is " SMBALERT_NI1->I2C1_SCL_F2H_SCP=-0.284";
   attribute ment_tsu302: string;
   attribute ment_tsu302 of DEF_ARCH : architecture is " SMBSUS_NI0->I2C0_SCL_F2H_SCP=-0.778";
   attribute ment_tsu303: string;
   attribute ment_tsu303 of DEF_ARCH : architecture is " SMBSUS_NI1->I2C1_SCL_F2H_SCP=-0.476";
   attribute ment_tsu304: string;
   attribute ment_tsu304 of DEF_ARCH : architecture is " SPI0_SDI_F2H_SCP->SPI0_CLK_IN=-0.010";
   attribute ment_tsu305: string;
   attribute ment_tsu305 of DEF_ARCH : architecture is " SPI1_SDI_F2H_SCP->SPI1_CLK_IN=-0.195";
   attribute ment_tco0: string;
   attribute ment_tco0 of DEF_ARCH : architecture is " CLK_BASE->CAN_RXBUS_MGPIO3A_H2F_A=3.441";
   attribute ment_tco1: string;
   attribute ment_tco1 of DEF_ARCH : architecture is " CLK_BASE->CAN_RXBUS_MGPIO3A_H2F_B=3.282";
   attribute ment_tco2: string;
   attribute ment_tco2 of DEF_ARCH : architecture is " CLK_BASE->CAN_TXBUS_MGPIO2A_H2F_A=3.471";
   attribute ment_tco3: string;
   attribute ment_tco3 of DEF_ARCH : architecture is " CLK_BASE->CAN_TXBUS_MGPIO2A_H2F_B=3.470";
   attribute ment_tco4: string;
   attribute ment_tco4 of DEF_ARCH : architecture is " CLK_BASE->CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT=3.711";
   attribute ment_tco5: string;
   attribute ment_tco5 of DEF_ARCH : architecture is " CLK_BASE->CAN_TX_EBL_MGPIO4A_H2F_A=3.345";
   attribute ment_tco6: string;
   attribute ment_tco6 of DEF_ARCH : architecture is " CLK_BASE->CAN_TX_EBL_MGPIO4A_H2F_B=3.542";
   attribute ment_tco7: string;
   attribute ment_tco7 of DEF_ARCH : architecture is " CLK_BASE->CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT=3.725";
   attribute ment_tco8: string;
   attribute ment_tco8 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[0]=3.882";
   attribute ment_tco9: string;
   attribute ment_tco9 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[10]=3.862";
   attribute ment_tco10: string;
   attribute ment_tco10 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[11]=3.866";
   attribute ment_tco11: string;
   attribute ment_tco11 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[12]=3.900";
   attribute ment_tco12: string;
   attribute ment_tco12 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[13]=3.906";
   attribute ment_tco13: string;
   attribute ment_tco13 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[14]=3.899";
   attribute ment_tco14: string;
   attribute ment_tco14 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[15]=3.914";
   attribute ment_tco15: string;
   attribute ment_tco15 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[16]=3.763";
   attribute ment_tco16: string;
   attribute ment_tco16 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[17]=3.745";
   attribute ment_tco17: string;
   attribute ment_tco17 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[18]=3.809";
   attribute ment_tco18: string;
   attribute ment_tco18 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[19]=3.771";
   attribute ment_tco19: string;
   attribute ment_tco19 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[1]=4.115";
   attribute ment_tco20: string;
   attribute ment_tco20 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[20]=3.744";
   attribute ment_tco21: string;
   attribute ment_tco21 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[21]=3.762";
   attribute ment_tco22: string;
   attribute ment_tco22 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[22]=3.784";
   attribute ment_tco23: string;
   attribute ment_tco23 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[23]=3.783";
   attribute ment_tco24: string;
   attribute ment_tco24 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[24]=3.867";
   attribute ment_tco25: string;
   attribute ment_tco25 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[25]=3.765";
   attribute ment_tco26: string;
   attribute ment_tco26 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[26]=3.820";
   attribute ment_tco27: string;
   attribute ment_tco27 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[27]=3.840";
   attribute ment_tco28: string;
   attribute ment_tco28 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[28]=3.774";
   attribute ment_tco29: string;
   attribute ment_tco29 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[29]=3.792";
   attribute ment_tco30: string;
   attribute ment_tco30 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[2]=3.885";
   attribute ment_tco31: string;
   attribute ment_tco31 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[30]=3.823";
   attribute ment_tco32: string;
   attribute ment_tco32 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[31]=3.835";
   attribute ment_tco33: string;
   attribute ment_tco33 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[3]=3.865";
   attribute ment_tco34: string;
   attribute ment_tco34 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[4]=3.894";
   attribute ment_tco35: string;
   attribute ment_tco35 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[5]=3.883";
   attribute ment_tco36: string;
   attribute ment_tco36 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[6]=3.886";
   attribute ment_tco37: string;
   attribute ment_tco37 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[7]=3.911";
   attribute ment_tco38: string;
   attribute ment_tco38 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[8]=3.909";
   attribute ment_tco39: string;
   attribute ment_tco39 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[9]=3.870";
   attribute ment_tco40: string;
   attribute ment_tco40 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_READYOUT=3.526";
   attribute ment_tco41: string;
   attribute ment_tco41 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RESP=3.323";
   attribute ment_tco42: string;
   attribute ment_tco42 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[0]=3.651";
   attribute ment_tco43: string;
   attribute ment_tco43 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[10]=3.584";
   attribute ment_tco44: string;
   attribute ment_tco44 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[11]=3.579";
   attribute ment_tco45: string;
   attribute ment_tco45 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[12]=3.598";
   attribute ment_tco46: string;
   attribute ment_tco46 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[13]=3.591";
   attribute ment_tco47: string;
   attribute ment_tco47 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[14]=3.593";
   attribute ment_tco48: string;
   attribute ment_tco48 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[15]=3.596";
   attribute ment_tco49: string;
   attribute ment_tco49 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[16]=3.430";
   attribute ment_tco50: string;
   attribute ment_tco50 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[17]=3.345";
   attribute ment_tco51: string;
   attribute ment_tco51 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[18]=3.422";
   attribute ment_tco52: string;
   attribute ment_tco52 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[19]=3.464";
   attribute ment_tco53: string;
   attribute ment_tco53 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[1]=3.587";
   attribute ment_tco54: string;
   attribute ment_tco54 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[20]=3.353";
   attribute ment_tco55: string;
   attribute ment_tco55 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[21]=3.363";
   attribute ment_tco56: string;
   attribute ment_tco56 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[22]=3.455";
   attribute ment_tco57: string;
   attribute ment_tco57 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[23]=3.437";
   attribute ment_tco58: string;
   attribute ment_tco58 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[24]=3.442";
   attribute ment_tco59: string;
   attribute ment_tco59 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[25]=3.385";
   attribute ment_tco60: string;
   attribute ment_tco60 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[26]=3.351";
   attribute ment_tco61: string;
   attribute ment_tco61 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[27]=3.473";
   attribute ment_tco62: string;
   attribute ment_tco62 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[28]=3.485";
   attribute ment_tco63: string;
   attribute ment_tco63 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[29]=3.351";
   attribute ment_tco64: string;
   attribute ment_tco64 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[2]=3.514";
   attribute ment_tco65: string;
   attribute ment_tco65 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[30]=3.385";
   attribute ment_tco66: string;
   attribute ment_tco66 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[31]=3.367";
   attribute ment_tco67: string;
   attribute ment_tco67 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[3]=3.556";
   attribute ment_tco68: string;
   attribute ment_tco68 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[4]=3.580";
   attribute ment_tco69: string;
   attribute ment_tco69 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[5]=3.586";
   attribute ment_tco70: string;
   attribute ment_tco70 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[6]=3.526";
   attribute ment_tco71: string;
   attribute ment_tco71 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[7]=3.539";
   attribute ment_tco72: string;
   attribute ment_tco72 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[8]=3.581";
   attribute ment_tco73: string;
   attribute ment_tco73 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RDATA[9]=3.590";
   attribute ment_tco74: string;
   attribute ment_tco74 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_READYOUT=3.112";
   attribute ment_tco75: string;
   attribute ment_tco75 of DEF_ARCH : architecture is " CLK_BASE->F_FM1_RESP=3.001";
   attribute ment_tco76: string;
   attribute ment_tco76 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[0]=2.959";
   attribute ment_tco77: string;
   attribute ment_tco77 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[10]=2.977";
   attribute ment_tco78: string;
   attribute ment_tco78 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[11]=2.934";
   attribute ment_tco79: string;
   attribute ment_tco79 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[12]=3.053";
   attribute ment_tco80: string;
   attribute ment_tco80 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[13]=2.855";
   attribute ment_tco81: string;
   attribute ment_tco81 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[14]=2.856";
   attribute ment_tco82: string;
   attribute ment_tco82 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[15]=2.899";
   attribute ment_tco83: string;
   attribute ment_tco83 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[16]=2.724";
   attribute ment_tco84: string;
   attribute ment_tco84 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[17]=2.927";
   attribute ment_tco85: string;
   attribute ment_tco85 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[18]=2.859";
   attribute ment_tco86: string;
   attribute ment_tco86 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[19]=2.899";
   attribute ment_tco87: string;
   attribute ment_tco87 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[1]=2.952";
   attribute ment_tco88: string;
   attribute ment_tco88 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[20]=2.912";
   attribute ment_tco89: string;
   attribute ment_tco89 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[21]=2.914";
   attribute ment_tco90: string;
   attribute ment_tco90 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[22]=2.914";
   attribute ment_tco91: string;
   attribute ment_tco91 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[23]=2.912";
   attribute ment_tco92: string;
   attribute ment_tco92 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[24]=2.907";
   attribute ment_tco93: string;
   attribute ment_tco93 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[25]=2.944";
   attribute ment_tco94: string;
   attribute ment_tco94 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[26]=2.886";
   attribute ment_tco95: string;
   attribute ment_tco95 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[27]=2.928";
   attribute ment_tco96: string;
   attribute ment_tco96 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[28]=2.913";
   attribute ment_tco97: string;
   attribute ment_tco97 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[29]=2.920";
   attribute ment_tco98: string;
   attribute ment_tco98 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[2]=2.892";
   attribute ment_tco99: string;
   attribute ment_tco99 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[30]=2.877";
   attribute ment_tco100: string;
   attribute ment_tco100 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[31]=3.001";
   attribute ment_tco101: string;
   attribute ment_tco101 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[3]=2.979";
   attribute ment_tco102: string;
   attribute ment_tco102 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[4]=2.903";
   attribute ment_tco103: string;
   attribute ment_tco103 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[5]=2.864";
   attribute ment_tco104: string;
   attribute ment_tco104 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[6]=2.866";
   attribute ment_tco105: string;
   attribute ment_tco105 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[7]=2.867";
   attribute ment_tco106: string;
   attribute ment_tco106 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[8]=2.940";
   attribute ment_tco107: string;
   attribute ment_tco107 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[9]=2.883";
   attribute ment_tco108: string;
   attribute ment_tco108 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_SEL=2.986";
   attribute ment_tco109: string;
   attribute ment_tco109 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_SIZE[0]=2.862";
   attribute ment_tco110: string;
   attribute ment_tco110 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_SIZE[1]=2.870";
   attribute ment_tco111: string;
   attribute ment_tco111 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_TRANS1=2.955";
   attribute ment_tco112: string;
   attribute ment_tco112 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[0]=2.844";
   attribute ment_tco113: string;
   attribute ment_tco113 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[10]=2.937";
   attribute ment_tco114: string;
   attribute ment_tco114 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[11]=2.912";
   attribute ment_tco115: string;
   attribute ment_tco115 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[12]=2.847";
   attribute ment_tco116: string;
   attribute ment_tco116 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[13]=3.009";
   attribute ment_tco117: string;
   attribute ment_tco117 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[14]=2.895";
   attribute ment_tco118: string;
   attribute ment_tco118 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[15]=2.908";
   attribute ment_tco119: string;
   attribute ment_tco119 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[16]=2.941";
   attribute ment_tco120: string;
   attribute ment_tco120 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[17]=2.941";
   attribute ment_tco121: string;
   attribute ment_tco121 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[18]=2.944";
   attribute ment_tco122: string;
   attribute ment_tco122 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[19]=2.859";
   attribute ment_tco123: string;
   attribute ment_tco123 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[1]=2.963";
   attribute ment_tco124: string;
   attribute ment_tco124 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[20]=2.895";
   attribute ment_tco125: string;
   attribute ment_tco125 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[21]=2.904";
   attribute ment_tco126: string;
   attribute ment_tco126 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[22]=2.928";
   attribute ment_tco127: string;
   attribute ment_tco127 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[23]=2.876";
   attribute ment_tco128: string;
   attribute ment_tco128 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[24]=2.884";
   attribute ment_tco129: string;
   attribute ment_tco129 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[25]=2.977";
   attribute ment_tco130: string;
   attribute ment_tco130 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[26]=2.928";
   attribute ment_tco131: string;
   attribute ment_tco131 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[27]=2.890";
   attribute ment_tco132: string;
   attribute ment_tco132 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[28]=2.854";
   attribute ment_tco133: string;
   attribute ment_tco133 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[29]=2.993";
   attribute ment_tco134: string;
   attribute ment_tco134 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[2]=2.860";
   attribute ment_tco135: string;
   attribute ment_tco135 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[30]=2.911";
   attribute ment_tco136: string;
   attribute ment_tco136 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[31]=2.905";
   attribute ment_tco137: string;
   attribute ment_tco137 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[3]=2.923";
   attribute ment_tco138: string;
   attribute ment_tco138 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[4]=2.907";
   attribute ment_tco139: string;
   attribute ment_tco139 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[5]=2.886";
   attribute ment_tco140: string;
   attribute ment_tco140 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[6]=2.879";
   attribute ment_tco141: string;
   attribute ment_tco141 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[7]=3.050";
   attribute ment_tco142: string;
   attribute ment_tco142 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[8]=2.996";
   attribute ment_tco143: string;
   attribute ment_tco143 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[9]=2.925";
   attribute ment_tco144: string;
   attribute ment_tco144 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WRITE=2.905";
   attribute ment_tco145: string;
   attribute ment_tco145 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[0]=2.786";
   attribute ment_tco146: string;
   attribute ment_tco146 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[10]=3.052";
   attribute ment_tco147: string;
   attribute ment_tco147 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[11]=2.757";
   attribute ment_tco148: string;
   attribute ment_tco148 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[12]=2.992";
   attribute ment_tco149: string;
   attribute ment_tco149 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[13]=2.802";
   attribute ment_tco150: string;
   attribute ment_tco150 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[14]=2.949";
   attribute ment_tco151: string;
   attribute ment_tco151 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[15]=2.746";
   attribute ment_tco152: string;
   attribute ment_tco152 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[16]=2.756";
   attribute ment_tco153: string;
   attribute ment_tco153 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[17]=2.771";
   attribute ment_tco154: string;
   attribute ment_tco154 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[18]=2.791";
   attribute ment_tco155: string;
   attribute ment_tco155 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[19]=2.868";
   attribute ment_tco156: string;
   attribute ment_tco156 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[1]=2.858";
   attribute ment_tco157: string;
   attribute ment_tco157 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[20]=2.891";
   attribute ment_tco158: string;
   attribute ment_tco158 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[21]=2.765";
   attribute ment_tco159: string;
   attribute ment_tco159 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[22]=2.760";
   attribute ment_tco160: string;
   attribute ment_tco160 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[23]=2.897";
   attribute ment_tco161: string;
   attribute ment_tco161 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[24]=2.717";
   attribute ment_tco162: string;
   attribute ment_tco162 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[25]=2.704";
   attribute ment_tco163: string;
   attribute ment_tco163 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[26]=2.693";
   attribute ment_tco164: string;
   attribute ment_tco164 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[27]=2.723";
   attribute ment_tco165: string;
   attribute ment_tco165 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[28]=2.711";
   attribute ment_tco166: string;
   attribute ment_tco166 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[29]=2.711";
   attribute ment_tco167: string;
   attribute ment_tco167 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[2]=2.858";
   attribute ment_tco168: string;
   attribute ment_tco168 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[30]=2.723";
   attribute ment_tco169: string;
   attribute ment_tco169 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[31]=2.728";
   attribute ment_tco170: string;
   attribute ment_tco170 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[3]=2.962";
   attribute ment_tco171: string;
   attribute ment_tco171 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[4]=2.891";
   attribute ment_tco172: string;
   attribute ment_tco172 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[5]=2.901";
   attribute ment_tco173: string;
   attribute ment_tco173 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[6]=2.876";
   attribute ment_tco174: string;
   attribute ment_tco174 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[7]=2.865";
   attribute ment_tco175: string;
   attribute ment_tco175 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[8]=2.931";
   attribute ment_tco176: string;
   attribute ment_tco176 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ADDR[9]=2.950";
   attribute ment_tco177: string;
   attribute ment_tco177 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_ENABLE=2.919";
   attribute ment_tco178: string;
   attribute ment_tco178 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_SEL=2.948";
   attribute ment_tco179: string;
   attribute ment_tco179 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[0]=2.781";
   attribute ment_tco180: string;
   attribute ment_tco180 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[10]=2.887";
   attribute ment_tco181: string;
   attribute ment_tco181 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[11]=2.867";
   attribute ment_tco182: string;
   attribute ment_tco182 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[12]=2.896";
   attribute ment_tco183: string;
   attribute ment_tco183 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[13]=2.890";
   attribute ment_tco184: string;
   attribute ment_tco184 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[14]=2.855";
   attribute ment_tco185: string;
   attribute ment_tco185 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[15]=2.864";
   attribute ment_tco186: string;
   attribute ment_tco186 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[16]=2.867";
   attribute ment_tco187: string;
   attribute ment_tco187 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[17]=2.844";
   attribute ment_tco188: string;
   attribute ment_tco188 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[18]=2.831";
   attribute ment_tco189: string;
   attribute ment_tco189 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[19]=2.849";
   attribute ment_tco190: string;
   attribute ment_tco190 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[1]=2.863";
   attribute ment_tco191: string;
   attribute ment_tco191 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[20]=2.804";
   attribute ment_tco192: string;
   attribute ment_tco192 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[21]=2.959";
   attribute ment_tco193: string;
   attribute ment_tco193 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[22]=2.943";
   attribute ment_tco194: string;
   attribute ment_tco194 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[23]=2.954";
   attribute ment_tco195: string;
   attribute ment_tco195 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[24]=2.935";
   attribute ment_tco196: string;
   attribute ment_tco196 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[25]=2.953";
   attribute ment_tco197: string;
   attribute ment_tco197 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[26]=2.799";
   attribute ment_tco198: string;
   attribute ment_tco198 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[27]=2.932";
   attribute ment_tco199: string;
   attribute ment_tco199 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[28]=2.828";
   attribute ment_tco200: string;
   attribute ment_tco200 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[29]=2.928";
   attribute ment_tco201: string;
   attribute ment_tco201 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[2]=2.929";
   attribute ment_tco202: string;
   attribute ment_tco202 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[30]=2.917";
   attribute ment_tco203: string;
   attribute ment_tco203 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[31]=2.961";
   attribute ment_tco204: string;
   attribute ment_tco204 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[3]=2.766";
   attribute ment_tco205: string;
   attribute ment_tco205 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[4]=2.831";
   attribute ment_tco206: string;
   attribute ment_tco206 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[5]=3.006";
   attribute ment_tco207: string;
   attribute ment_tco207 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[6]=2.864";
   attribute ment_tco208: string;
   attribute ment_tco208 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[7]=2.942";
   attribute ment_tco209: string;
   attribute ment_tco209 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[8]=2.904";
   attribute ment_tco210: string;
   attribute ment_tco210 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WDATA[9]=2.844";
   attribute ment_tco211: string;
   attribute ment_tco211 of DEF_ARCH : architecture is " CLK_BASE->F_HM1_WRITE=3.150";
   attribute ment_tco212: string;
   attribute ment_tco212 of DEF_ARCH : architecture is " CLK_BASE->H2FCALIB=3.130";
   attribute ment_tco213: string;
   attribute ment_tco213 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SCL_MGPIO31B_H2F_B=3.603";
   attribute ment_tco214: string;
   attribute ment_tco214 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SCL_USBC_DATA1_MGPIO31B_OE=2.746";
   attribute ment_tco215: string;
   attribute ment_tco215 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SDA_MGPIO30B_H2F_A=3.520";
   attribute ment_tco216: string;
   attribute ment_tco216 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SDA_MGPIO30B_H2F_B=3.581";
   attribute ment_tco217: string;
   attribute ment_tco217 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SDA_USBC_DATA0_MGPIO30B_OE=2.887";
   attribute ment_tco218: string;
   attribute ment_tco218 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SCL_MGPIO1A_H2F_B=3.320";
   attribute ment_tco219: string;
   attribute ment_tco219 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SCL_USBA_DATA4_MGPIO1A_OE=3.266";
   attribute ment_tco220: string;
   attribute ment_tco220 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SDA_MGPIO0A_H2F_A=3.613";
   attribute ment_tco221: string;
   attribute ment_tco221 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SDA_MGPIO0A_H2F_B=3.522";
   attribute ment_tco222: string;
   attribute ment_tco222 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SDA_USBA_DATA3_MGPIO0A_OE=3.166";
   attribute ment_tco223: string;
   attribute ment_tco223 of DEF_ARCH : architecture is " CLK_BASE->MGPIO0B_OE=2.062";
   attribute ment_tco224: string;
   attribute ment_tco224 of DEF_ARCH : architecture is " CLK_BASE->MGPIO0B_OUT=1.940";
   attribute ment_tco225: string;
   attribute ment_tco225 of DEF_ARCH : architecture is " CLK_BASE->MGPIO10B_OE=2.578";
   attribute ment_tco226: string;
   attribute ment_tco226 of DEF_ARCH : architecture is " CLK_BASE->MGPIO10B_OUT=2.432";
   attribute ment_tco227: string;
   attribute ment_tco227 of DEF_ARCH : architecture is " CLK_BASE->MGPIO1B_OE=1.997";
   attribute ment_tco228: string;
   attribute ment_tco228 of DEF_ARCH : architecture is " CLK_BASE->MGPIO1B_OUT=1.993";
   attribute ment_tco229: string;
   attribute ment_tco229 of DEF_ARCH : architecture is " CLK_BASE->MGPIO25A_OE=2.105";
   attribute ment_tco230: string;
   attribute ment_tco230 of DEF_ARCH : architecture is " CLK_BASE->MGPIO25A_OUT=2.516";
   attribute ment_tco231: string;
   attribute ment_tco231 of DEF_ARCH : architecture is " CLK_BASE->MGPIO26A_OE=2.099";
   attribute ment_tco232: string;
   attribute ment_tco232 of DEF_ARCH : architecture is " CLK_BASE->MGPIO26A_OUT=2.174";
   attribute ment_tco233: string;
   attribute ment_tco233 of DEF_ARCH : architecture is " CLK_BASE->MGPIO27A_OE=3.236";
   attribute ment_tco234: string;
   attribute ment_tco234 of DEF_ARCH : architecture is " CLK_BASE->MGPIO27A_OUT=3.473";
   attribute ment_tco235: string;
   attribute ment_tco235 of DEF_ARCH : architecture is " CLK_BASE->MGPIO28A_OE=3.587";
   attribute ment_tco236: string;
   attribute ment_tco236 of DEF_ARCH : architecture is " CLK_BASE->MGPIO28A_OUT=3.281";
   attribute ment_tco237: string;
   attribute ment_tco237 of DEF_ARCH : architecture is " CLK_BASE->MGPIO29A_OE=2.035";
   attribute ment_tco238: string;
   attribute ment_tco238 of DEF_ARCH : architecture is " CLK_BASE->MGPIO29A_OUT=1.973";
   attribute ment_tco239: string;
   attribute ment_tco239 of DEF_ARCH : architecture is " CLK_BASE->MGPIO2B_OE=2.100";
   attribute ment_tco240: string;
   attribute ment_tco240 of DEF_ARCH : architecture is " CLK_BASE->MGPIO2B_OUT=2.055";
   attribute ment_tco241: string;
   attribute ment_tco241 of DEF_ARCH : architecture is " CLK_BASE->MGPIO30A_OE=2.036";
   attribute ment_tco242: string;
   attribute ment_tco242 of DEF_ARCH : architecture is " CLK_BASE->MGPIO30A_OUT=2.036";
   attribute ment_tco243: string;
   attribute ment_tco243 of DEF_ARCH : architecture is " CLK_BASE->MGPIO31A_OE=1.935";
   attribute ment_tco244: string;
   attribute ment_tco244 of DEF_ARCH : architecture is " CLK_BASE->MGPIO31A_OUT=1.912";
   attribute ment_tco245: string;
   attribute ment_tco245 of DEF_ARCH : architecture is " CLK_BASE->MGPIO3B_OE=2.153";
   attribute ment_tco246: string;
   attribute ment_tco246 of DEF_ARCH : architecture is " CLK_BASE->MGPIO3B_OUT=2.294";
   attribute ment_tco247: string;
   attribute ment_tco247 of DEF_ARCH : architecture is " CLK_BASE->MGPIO4B_OE=2.243";
   attribute ment_tco248: string;
   attribute ment_tco248 of DEF_ARCH : architecture is " CLK_BASE->MGPIO4B_OUT=2.615";
   attribute ment_tco249: string;
   attribute ment_tco249 of DEF_ARCH : architecture is " CLK_BASE->MGPIO5B_OE=2.498";
   attribute ment_tco250: string;
   attribute ment_tco250 of DEF_ARCH : architecture is " CLK_BASE->MGPIO5B_OUT=2.841";
   attribute ment_tco251: string;
   attribute ment_tco251 of DEF_ARCH : architecture is " CLK_BASE->MGPIO6B_OE=2.779";
   attribute ment_tco252: string;
   attribute ment_tco252 of DEF_ARCH : architecture is " CLK_BASE->MGPIO6B_OUT=2.489";
   attribute ment_tco253: string;
   attribute ment_tco253 of DEF_ARCH : architecture is " CLK_BASE->MGPIO7B_OE=2.391";
   attribute ment_tco254: string;
   attribute ment_tco254 of DEF_ARCH : architecture is " CLK_BASE->MGPIO7B_OUT=2.379";
   attribute ment_tco255: string;
   attribute ment_tco255 of DEF_ARCH : architecture is " CLK_BASE->MGPIO8B_OE=2.273";
   attribute ment_tco256: string;
   attribute ment_tco256 of DEF_ARCH : architecture is " CLK_BASE->MGPIO8B_OUT=2.441";
   attribute ment_tco257: string;
   attribute ment_tco257 of DEF_ARCH : architecture is " CLK_BASE->MGPIO9B_OE=2.273";
   attribute ment_tco258: string;
   attribute ment_tco258 of DEF_ARCH : architecture is " CLK_BASE->MGPIO9B_OUT=2.474";
   attribute ment_tco259: string;
   attribute ment_tco259 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_CTS_MGPIO19B_H2F_A=3.375";
   attribute ment_tco260: string;
   attribute ment_tco260 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_CTS_MGPIO19B_H2F_B=3.377";
   attribute ment_tco261: string;
   attribute ment_tco261 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DCD_MGPIO22B_H2F_A=3.445";
   attribute ment_tco262: string;
   attribute ment_tco262 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DCD_MGPIO22B_H2F_B=3.518";
   attribute ment_tco263: string;
   attribute ment_tco263 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DSR_MGPIO20B_H2F_A=3.411";
   attribute ment_tco264: string;
   attribute ment_tco264 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DSR_MGPIO20B_H2F_B=3.655";
   attribute ment_tco265: string;
   attribute ment_tco265 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DTR_MGPIO18B_H2F_A=3.270";
   attribute ment_tco266: string;
   attribute ment_tco266 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DTR_MGPIO18B_H2F_B=3.480";
   attribute ment_tco267: string;
   attribute ment_tco267 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT=2.658";
   attribute ment_tco268: string;
   attribute ment_tco268 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RI_MGPIO21B_H2F_A=3.523";
   attribute ment_tco269: string;
   attribute ment_tco269 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RI_MGPIO21B_H2F_B=3.764";
   attribute ment_tco270: string;
   attribute ment_tco270 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RTS_MGPIO17B_H2F_A=3.587";
   attribute ment_tco271: string;
   attribute ment_tco271 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RTS_MGPIO17B_H2F_B=3.320";
   attribute ment_tco272: string;
   attribute ment_tco272 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT=2.689";
   attribute ment_tco273: string;
   attribute ment_tco273 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RXD_MGPIO28B_H2F_A=3.714";
   attribute ment_tco274: string;
   attribute ment_tco274 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RXD_MGPIO28B_H2F_B=3.566";
   attribute ment_tco275: string;
   attribute ment_tco275 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_SCK_MGPIO29B_H2F_A=3.380";
   attribute ment_tco276: string;
   attribute ment_tco276 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_SCK_MGPIO29B_H2F_B=3.646";
   attribute ment_tco277: string;
   attribute ment_tco277 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_SCK_USBC_NXT_MGPIO29B_OE=3.584";
   attribute ment_tco278: string;
   attribute ment_tco278 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_SCK_USBC_NXT_MGPIO29B_OUT=2.765";
   attribute ment_tco279: string;
   attribute ment_tco279 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_TXD_MGPIO27B_H2F_A=3.879";
   attribute ment_tco280: string;
   attribute ment_tco280 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_TXD_MGPIO27B_H2F_B=3.839";
   attribute ment_tco281: string;
   attribute ment_tco281 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_TXD_USBC_DIR_MGPIO27B_OE=3.162";
   attribute ment_tco282: string;
   attribute ment_tco282 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_TXD_USBC_DIR_MGPIO27B_OUT=3.243";
   attribute ment_tco283: string;
   attribute ment_tco283 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_DTR_MGPIO12B_H2F_A=3.713";
   attribute ment_tco284: string;
   attribute ment_tco284 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_DTR_MGPIO12B_OUT=3.609";
   attribute ment_tco285: string;
   attribute ment_tco285 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RTS_MGPIO11B_H2F_A=3.534";
   attribute ment_tco286: string;
   attribute ment_tco286 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RTS_MGPIO11B_H2F_B=3.508";
   attribute ment_tco287: string;
   attribute ment_tco287 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RTS_MGPIO11B_OUT=3.762";
   attribute ment_tco288: string;
   attribute ment_tco288 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RXD_MGPIO26B_H2F_A=3.653";
   attribute ment_tco289: string;
   attribute ment_tco289 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RXD_MGPIO26B_H2F_B=3.470";
   attribute ment_tco290: string;
   attribute ment_tco290 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_SCK_MGPIO25B_H2F_A=3.515";
   attribute ment_tco291: string;
   attribute ment_tco291 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_SCK_MGPIO25B_H2F_B=3.969";
   attribute ment_tco292: string;
   attribute ment_tco292 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_SCK_USBC_DATA4_MGPIO25B_OE=4.211";
   attribute ment_tco293: string;
   attribute ment_tco293 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT=3.481";
   attribute ment_tco294: string;
   attribute ment_tco294 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_TXD_MGPIO24B_H2F_A=3.506";
   attribute ment_tco295: string;
   attribute ment_tco295 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_TXD_MGPIO24B_H2F_B=3.598";
   attribute ment_tco296: string;
   attribute ment_tco296 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_TXD_USBC_DATA2_MGPIO24B_OE=4.053";
   attribute ment_tco297: string;
   attribute ment_tco297 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT=3.955";
   attribute ment_tco298: string;
   attribute ment_tco298 of DEF_ARCH : architecture is " CLK_BASE->RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE=4.174";
   attribute ment_tco299: string;
   attribute ment_tco299 of DEF_ARCH : architecture is " CLK_BASE->RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT=3.528";
   attribute ment_tco300: string;
   attribute ment_tco300 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDI_MGPIO5A_H2F_A=3.447";
   attribute ment_tco301: string;
   attribute ment_tco301 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDI_MGPIO5A_H2F_B=3.758";
   attribute ment_tco302: string;
   attribute ment_tco302 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDO_MGPIO6A_H2F_A=3.966";
   attribute ment_tco303: string;
   attribute ment_tco303 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDO_MGPIO6A_H2F_B=3.813";
   attribute ment_tco304: string;
   attribute ment_tco304 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDO_USBA_STP_MGPIO6A_OE=4.755";
   attribute ment_tco305: string;
   attribute ment_tco305 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDO_USBA_STP_MGPIO6A_OUT=4.301";
   attribute ment_tco306: string;
   attribute ment_tco306 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS0_MGPIO7A_H2F_A=3.421";
   attribute ment_tco307: string;
   attribute ment_tco307 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS0_MGPIO7A_H2F_B=3.641";
   attribute ment_tco308: string;
   attribute ment_tco308 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS1_MGPIO8A_H2F_A=3.297";
   attribute ment_tco309: string;
   attribute ment_tco309 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS1_MGPIO8A_H2F_B=3.620";
   attribute ment_tco310: string;
   attribute ment_tco310 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS2_MGPIO9A_H2F_A=3.530";
   attribute ment_tco311: string;
   attribute ment_tco311 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS2_MGPIO9A_H2F_B=3.596";
   attribute ment_tco312: string;
   attribute ment_tco312 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS3_MGPIO10A_H2F_A=3.638";
   attribute ment_tco313: string;
   attribute ment_tco313 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS3_MGPIO10A_H2F_B=3.577";
   attribute ment_tco314: string;
   attribute ment_tco314 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS4_MGPIO19A_H2F_A=3.374";
   attribute ment_tco315: string;
   attribute ment_tco315 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS5_MGPIO20A_H2F_A=3.470";
   attribute ment_tco316: string;
   attribute ment_tco316 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS6_MGPIO21A_H2F_A=3.452";
   attribute ment_tco317: string;
   attribute ment_tco317 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS7_MGPIO22A_H2F_A=3.426";
   attribute ment_tco318: string;
   attribute ment_tco318 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDI_MGPIO11A_H2F_A=3.509";
   attribute ment_tco319: string;
   attribute ment_tco319 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDI_MGPIO11A_H2F_B=3.471";
   attribute ment_tco320: string;
   attribute ment_tco320 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDO_MGPIO12A_H2F_A=3.850";
   attribute ment_tco321: string;
   attribute ment_tco321 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDO_MGPIO12A_H2F_B=3.804";
   attribute ment_tco322: string;
   attribute ment_tco322 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDO_MGPIO12A_OE=6.223";
   attribute ment_tco323: string;
   attribute ment_tco323 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDO_MGPIO12A_OUT=5.639";
   attribute ment_tco324: string;
   attribute ment_tco324 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS0_MGPIO13A_H2F_A=3.818";
   attribute ment_tco325: string;
   attribute ment_tco325 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS0_MGPIO13A_H2F_B=3.556";
   attribute ment_tco326: string;
   attribute ment_tco326 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS1_MGPIO14A_H2F_A=3.636";
   attribute ment_tco327: string;
   attribute ment_tco327 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS1_MGPIO14A_H2F_B=3.405";
   attribute ment_tco328: string;
   attribute ment_tco328 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS2_MGPIO15A_H2F_A=3.448";
   attribute ment_tco329: string;
   attribute ment_tco329 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS2_MGPIO15A_H2F_B=3.405";
   attribute ment_tco330: string;
   attribute ment_tco330 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS3_MGPIO16A_H2F_A=3.600";
   attribute ment_tco331: string;
   attribute ment_tco331 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS3_MGPIO16A_H2F_B=3.574";
   attribute ment_tco332: string;
   attribute ment_tco332 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS4_MGPIO17A_H2F_A=3.522";
   attribute ment_tco333: string;
   attribute ment_tco333 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS5_MGPIO18A_H2F_A=3.312";
   attribute ment_tco334: string;
   attribute ment_tco334 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS6_MGPIO23A_H2F_A=3.527";
   attribute ment_tco335: string;
   attribute ment_tco335 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS7_MGPIO24A_H2F_A=3.489";
   attribute ment_tco336: string;
   attribute ment_tco336 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PRDATA[0]=8.740";
   attribute ment_tco337: string;
   attribute ment_tco337 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PRDATA[10]=4.987";
   attribute ment_tco338: string;
   attribute ment_tco338 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PRDATA[11]=5.034";
   attribute ment_tco339: string;
   attribute ment_tco339 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PRDATA[12]=4.958";
   attribute ment_tco340: string;
   attribute ment_tco340 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PRDATA[13]=4.775";
   attribute ment_tco341: string;
   attribute ment_tco341 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PRDATA[14]=4.842";
   attribute ment_tco342: string;
   attribute ment_tco342 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PRDATA[15]=4.923";
   attribute ment_tco343: string;
   attribute ment_tco343 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PRDATA[1]=8.660";
   attribute ment_tco344: string;
   attribute ment_tco344 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PRDATA[2]=8.366";
   attribute ment_tco345: string;
   attribute ment_tco345 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PRDATA[3]=8.960";
   attribute ment_tco346: string;
   attribute ment_tco346 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PRDATA[4]=4.776";
   attribute ment_tco347: string;
   attribute ment_tco347 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PRDATA[5]=5.038";
   attribute ment_tco348: string;
   attribute ment_tco348 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PRDATA[6]=4.788";
   attribute ment_tco349: string;
   attribute ment_tco349 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PRDATA[7]=4.891";
   attribute ment_tco350: string;
   attribute ment_tco350 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PRDATA[8]=4.954";
   attribute ment_tco351: string;
   attribute ment_tco351 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PRDATA[9]=4.916";
   attribute ment_tco352: string;
   attribute ment_tco352 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PREADY=5.147";
   attribute ment_tco353: string;
   attribute ment_tco353 of DEF_ARCH : architecture is " CLK_MDDR_APB->MDDR_FABRIC_PSLVERR=4.262";
   attribute black_box_pad : string;
   attribute black_box_pad of DEF_ARCH : architecture is "";

begin

end DEF_ARCH;
