../../../rtl/ram_mux.vhd