../../../rtl/orca.vhd