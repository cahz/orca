../../../rtl/instruction_fetch.vhd