../../../rtl/sys_call.vhd