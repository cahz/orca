../../../rtl/microsemi_wrapper.vhd