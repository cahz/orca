../../rtl/utils.vhd