../../../rtl/branch_unit.vhd