../../../rtl/alu.vhd