../../../rtl/bram_microsemi.vhd