//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Fri Jun 16 12:00:37 2017
// Version: v11.7 SP3 11.7.3.8
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// tb
module tb(
);

//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   RESET_GEN_0_RESET;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire   GND_net;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign GND_net = 1'b0;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------RESET_GEN   -   Actel:Simulation:RESET_GEN:1.0.1
RESET_GEN #( 
        .DELAY       ( 500 ),
        .LOGIC_LEVEL ( 0 ) )
RESET_GEN_0(
        // Outputs
        .RESET ( RESET_GEN_0_RESET ) 
        );

//--------Top_Fabric_Master
Top_Fabric_Master Top_Fabric_Master_0(
        // Inputs
        .DEVRST_N ( RESET_GEN_0_RESET ),
        .RX       ( GND_net ),
        // Outputs
        .TX       (  ) 
        );


endmodule
