../../idram.vhd