../../rtl/orca.vhd