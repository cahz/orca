../../utils.vhd