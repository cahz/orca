../../edge_extender.vhd