../../../rtl/utils.vhd