../../../rtl/execute.vhd