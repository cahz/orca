../../../rtl/load_store_unit.vhd