../../rtl/axi_master.vhd