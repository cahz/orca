../../constants_pkg.vhd