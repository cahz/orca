../../../rtl/cache_xilinx.vhd