../../../rtl/register_file.vhd