../../components.vhd