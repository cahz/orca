../../rtl/constants_pkg.vhd