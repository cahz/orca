../../rtl/components.vhd