../../rtl/lve_top.vhd