../../../rtl/decode.vhd